library ieee;
use ieee.std_logic_1164.all;

library std;
use std.pkg_ram.all;

library bre;
use bre.pkg_bre.all;

entity top is
	Port (
		clk_i    :  in std_logic;
		rst_i    :  in std_logic;
		query_i  :  in query_in_array_type;
		result_o : out std_logic_vector(157 downto 0);
		mem_i    :  in std_logic_vector(200 downto 0);
		meme_i   :  in std_logic_vector(5 downto 0)
	);
end top;

architecture behavioural of top is
	signal sig_fnc_RTD	: std_logic_vector(2799 downto 0);
	signal sig_ram_VERS	: std_logic_vector(4 downto 0);
	signal sig_fnc_OWN	: std_logic_vector(1188 downto 0);
	signal sig_ram_APP	: std_logic_vector(44 downto 0);
	signal sig_fnc_DATE	: std_logic_vector(99 downto 0);
	signal sig_ram_MKTA	: std_logic_vector(31 downto 0);
	signal sig_ram_MKTB	: std_logic_vector(31 downto 0);
	signal sig_ram_CABIN	: std_logic_vector(7 downto 0);
	signal sig_ram_BKG	: std_logic_vector(25 downto 0);
begin

fnc_RTD0 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000000000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(0)
);
fnc_RTD1 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000000001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1)
);
fnc_RTD2 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000000010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2)
);
fnc_RTD3 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000000011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(3)
);
fnc_RTD4 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000000100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(4)
);
fnc_RTD5 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000000101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(5)
);
fnc_RTD6 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000000110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(6)
);
fnc_RTD7 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000000111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(7)
);
fnc_RTD8 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000001000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(8)
);
fnc_RTD9 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000001001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(9)
);
fnc_RTD10 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000001010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(10)
);
fnc_RTD11 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000001011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(11)
);
fnc_RTD12 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000001100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(12)
);
fnc_RTD13 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000001101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(13)
);
fnc_RTD14 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000001110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(14)
);
fnc_RTD15 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000001111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(15)
);
fnc_RTD16 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000010000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(16)
);
fnc_RTD17 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000010001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(17)
);
fnc_RTD18 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000010010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(18)
);
fnc_RTD19 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000010011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(19)
);
fnc_RTD20 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000010100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(20)
);
fnc_RTD21 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000010101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(21)
);
fnc_RTD22 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000010110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(22)
);
fnc_RTD23 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000010111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(23)
);
fnc_RTD24 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000011000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(24)
);
fnc_RTD25 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000011001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(25)
);
fnc_RTD26 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000011010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(26)
);
fnc_RTD27 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000011011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(27)
);
fnc_RTD28 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000011100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(28)
);
fnc_RTD29 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000011101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(29)
);
fnc_RTD30 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000011110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(30)
);
fnc_RTD31 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000011111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(31)
);
fnc_RTD32 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000100000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(32)
);
fnc_RTD33 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000100001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(33)
);
fnc_RTD34 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000100010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(34)
);
fnc_RTD35 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000100011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(35)
);
fnc_RTD36 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000100100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(36)
);
fnc_RTD37 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000100101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(37)
);
fnc_RTD38 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000100110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(38)
);
fnc_RTD39 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000100111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(39)
);
fnc_RTD40 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000101000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(40)
);
fnc_RTD41 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000101001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(41)
);
fnc_RTD42 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000101010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(42)
);
fnc_RTD43 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000101011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(43)
);
fnc_RTD44 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000101100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(44)
);
fnc_RTD45 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000101101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(45)
);
fnc_RTD46 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000101110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(46)
);
fnc_RTD47 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000101111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(47)
);
fnc_RTD48 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000110000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(48)
);
fnc_RTD49 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000110001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(49)
);
fnc_RTD50 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000110010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(50)
);
fnc_RTD51 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000110011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(51)
);
fnc_RTD52 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000110100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(52)
);
fnc_RTD53 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000110101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(53)
);
fnc_RTD54 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000110110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(54)
);
fnc_RTD55 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000110111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(55)
);
fnc_RTD56 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000111000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(56)
);
fnc_RTD57 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000111001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(57)
);
fnc_RTD58 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000111010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(58)
);
fnc_RTD59 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000111011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(59)
);
fnc_RTD60 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000111100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(60)
);
fnc_RTD61 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000111101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(61)
);
fnc_RTD62 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000111110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(62)
);
fnc_RTD63 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000111111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(63)
);
fnc_RTD64 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001000000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(64)
);
fnc_RTD65 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001000001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(65)
);
fnc_RTD66 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001000010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(66)
);
fnc_RTD67 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001000011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(67)
);
fnc_RTD68 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001000100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(68)
);
fnc_RTD69 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001000101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(69)
);
fnc_RTD70 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001000110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(70)
);
fnc_RTD71 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001000111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(71)
);
fnc_RTD72 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001001000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(72)
);
fnc_RTD73 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001001001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(73)
);
fnc_RTD74 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001001010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(74)
);
fnc_RTD75 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001001011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(75)
);
fnc_RTD76 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001001100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(76)
);
fnc_RTD77 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001001101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(77)
);
fnc_RTD78 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001001110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(78)
);
fnc_RTD79 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001001111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(79)
);
fnc_RTD80 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001010000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(80)
);
fnc_RTD81 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001010001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(81)
);
fnc_RTD82 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001010010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(82)
);
fnc_RTD83 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001010011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(83)
);
fnc_RTD84 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001010100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(84)
);
fnc_RTD85 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001010101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(85)
);
fnc_RTD86 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001010110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(86)
);
fnc_RTD87 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001010111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(87)
);
fnc_RTD88 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001011000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(88)
);
fnc_RTD89 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001011001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(89)
);
fnc_RTD90 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001011010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(90)
);
fnc_RTD91 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001011011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(91)
);
fnc_RTD92 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001011100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(92)
);
fnc_RTD93 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001011101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(93)
);
fnc_RTD94 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001011110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(94)
);
fnc_RTD95 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001011111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(95)
);
fnc_RTD96 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001100000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(96)
);
fnc_RTD97 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001100001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(97)
);
fnc_RTD98 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001100010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(98)
);
fnc_RTD99 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001100011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(99)
);
fnc_RTD100 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001100100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(100)
);
fnc_RTD101 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001100101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(101)
);
fnc_RTD102 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001100110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(102)
);
fnc_RTD103 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001100111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(103)
);
fnc_RTD104 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001101000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(104)
);
fnc_RTD105 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001101001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(105)
);
fnc_RTD106 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001101010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(106)
);
fnc_RTD107 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001101011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(107)
);
fnc_RTD108 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001101100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(108)
);
fnc_RTD109 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001101101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(109)
);
fnc_RTD110 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001101110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(110)
);
fnc_RTD111 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001101111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(111)
);
fnc_RTD112 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001110000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(112)
);
fnc_RTD113 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001110001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(113)
);
fnc_RTD114 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001110010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(114)
);
fnc_RTD115 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001110011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(115)
);
fnc_RTD116 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001110100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(116)
);
fnc_RTD117 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001110101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(117)
);
fnc_RTD118 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001110110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(118)
);
fnc_RTD119 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001110111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(119)
);
fnc_RTD120 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001111000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(120)
);
fnc_RTD121 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001111001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(121)
);
fnc_RTD122 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001111010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(122)
);
fnc_RTD123 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001111011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(123)
);
fnc_RTD124 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001111100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(124)
);
fnc_RTD125 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001111101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(125)
);
fnc_RTD126 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001111110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(126)
);
fnc_RTD127 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001111111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(127)
);
fnc_RTD128 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010000000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(128)
);
fnc_RTD129 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010000001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(129)
);
fnc_RTD130 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010000010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(130)
);
fnc_RTD131 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010000011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(131)
);
fnc_RTD132 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010000100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(132)
);
fnc_RTD133 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010000101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(133)
);
fnc_RTD134 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010000110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(134)
);
fnc_RTD135 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010000111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(135)
);
fnc_RTD136 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010001000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(136)
);
fnc_RTD137 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010001001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(137)
);
fnc_RTD138 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010001010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(138)
);
fnc_RTD139 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010001011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(139)
);
fnc_RTD140 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010001100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(140)
);
fnc_RTD141 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010001101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(141)
);
fnc_RTD142 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010001110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(142)
);
fnc_RTD143 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010001111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(143)
);
fnc_RTD144 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010010000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(144)
);
fnc_RTD145 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010010001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(145)
);
fnc_RTD146 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010010010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(146)
);
fnc_RTD147 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010010011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(147)
);
fnc_RTD148 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010010100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(148)
);
fnc_RTD149 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010010101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(149)
);
fnc_RTD150 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010010110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(150)
);
fnc_RTD151 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010010111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(151)
);
fnc_RTD152 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010011000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(152)
);
fnc_RTD153 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010011001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(153)
);
fnc_RTD154 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010011010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(154)
);
fnc_RTD155 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010011011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(155)
);
fnc_RTD156 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010011100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(156)
);
fnc_RTD157 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010011101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(157)
);
fnc_RTD158 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010011110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(158)
);
fnc_RTD159 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010011111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(159)
);
fnc_RTD160 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010100000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(160)
);
fnc_RTD161 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010100001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(161)
);
fnc_RTD162 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010100010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(162)
);
fnc_RTD163 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010100011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(163)
);
fnc_RTD164 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010100100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(164)
);
fnc_RTD165 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010100101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(165)
);
fnc_RTD166 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010100110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(166)
);
fnc_RTD167 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010100111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(167)
);
fnc_RTD168 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010101000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(168)
);
fnc_RTD169 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010101001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(169)
);
fnc_RTD170 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010101010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(170)
);
fnc_RTD171 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010101011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(171)
);
fnc_RTD172 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010101100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(172)
);
fnc_RTD173 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010101101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(173)
);
fnc_RTD174 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010101110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(174)
);
fnc_RTD175 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010101111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(175)
);
fnc_RTD176 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010110000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(176)
);
fnc_RTD177 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010110001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(177)
);
fnc_RTD178 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010110010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(178)
);
fnc_RTD179 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010110011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(179)
);
fnc_RTD180 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010110100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(180)
);
fnc_RTD181 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010110101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(181)
);
fnc_RTD182 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010110110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(182)
);
fnc_RTD183 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010110111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(183)
);
fnc_RTD184 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010111000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(184)
);
fnc_RTD185 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010111001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(185)
);
fnc_RTD186 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010111010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(186)
);
fnc_RTD187 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010111011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(187)
);
fnc_RTD188 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010111100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(188)
);
fnc_RTD189 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010111101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(189)
);
fnc_RTD190 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010111110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(190)
);
fnc_RTD191 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010111111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(191)
);
fnc_RTD192 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011000000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(192)
);
fnc_RTD193 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011000001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(193)
);
fnc_RTD194 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011000010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(194)
);
fnc_RTD195 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011000011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(195)
);
fnc_RTD196 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011000100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(196)
);
fnc_RTD197 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011000101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(197)
);
fnc_RTD198 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011000110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(198)
);
fnc_RTD199 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011000111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(199)
);
fnc_RTD200 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011001000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(200)
);
fnc_RTD201 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011001001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(201)
);
fnc_RTD202 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011001010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(202)
);
fnc_RTD203 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011001011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(203)
);
fnc_RTD204 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011001100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(204)
);
fnc_RTD205 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011001101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(205)
);
fnc_RTD206 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011001110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(206)
);
fnc_RTD207 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011001111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(207)
);
fnc_RTD208 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011010000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(208)
);
fnc_RTD209 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011010001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(209)
);
fnc_RTD210 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011010010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(210)
);
fnc_RTD211 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011010011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(211)
);
fnc_RTD212 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011010100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(212)
);
fnc_RTD213 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011010101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(213)
);
fnc_RTD214 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011010110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(214)
);
fnc_RTD215 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011010111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(215)
);
fnc_RTD216 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011011000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(216)
);
fnc_RTD217 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011011001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(217)
);
fnc_RTD218 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011011010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(218)
);
fnc_RTD219 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011011011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(219)
);
fnc_RTD220 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011011100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(220)
);
fnc_RTD221 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011011101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(221)
);
fnc_RTD222 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011011110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(222)
);
fnc_RTD223 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011011111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(223)
);
fnc_RTD224 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011100000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(224)
);
fnc_RTD225 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011100001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(225)
);
fnc_RTD226 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011100010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(226)
);
fnc_RTD227 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011100011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(227)
);
fnc_RTD228 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011100100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(228)
);
fnc_RTD229 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011100101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(229)
);
fnc_RTD230 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011100110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(230)
);
fnc_RTD231 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011100111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(231)
);
fnc_RTD232 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011101000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(232)
);
fnc_RTD233 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011101001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(233)
);
fnc_RTD234 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011101010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(234)
);
fnc_RTD235 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011101011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(235)
);
fnc_RTD236 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011101100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(236)
);
fnc_RTD237 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011101101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(237)
);
fnc_RTD238 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011101110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(238)
);
fnc_RTD239 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011101111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(239)
);
fnc_RTD240 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011110000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(240)
);
fnc_RTD241 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011110001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(241)
);
fnc_RTD242 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011110010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(242)
);
fnc_RTD243 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011110011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(243)
);
fnc_RTD244 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011110100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(244)
);
fnc_RTD245 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011110101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(245)
);
fnc_RTD246 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011110110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(246)
);
fnc_RTD247 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011110111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(247)
);
fnc_RTD248 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011111000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(248)
);
fnc_RTD249 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011111001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(249)
);
fnc_RTD250 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011111010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(250)
);
fnc_RTD251 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011111011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(251)
);
fnc_RTD252 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011111100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(252)
);
fnc_RTD253 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011111101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(253)
);
fnc_RTD254 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011111110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(254)
);
fnc_RTD255 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011111111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(255)
);
fnc_RTD256 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100000000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(256)
);
fnc_RTD257 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100000001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(257)
);
fnc_RTD258 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100000010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(258)
);
fnc_RTD259 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100000011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(259)
);
fnc_RTD260 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100000100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(260)
);
fnc_RTD261 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100000101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(261)
);
fnc_RTD262 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100000110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(262)
);
fnc_RTD263 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100000111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(263)
);
fnc_RTD264 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100001000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(264)
);
fnc_RTD265 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100001001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(265)
);
fnc_RTD266 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100001010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(266)
);
fnc_RTD267 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100001011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(267)
);
fnc_RTD268 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100001100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(268)
);
fnc_RTD269 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100001101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(269)
);
fnc_RTD270 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100001110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(270)
);
fnc_RTD271 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100001111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(271)
);
fnc_RTD272 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100010000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(272)
);
fnc_RTD273 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100010001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(273)
);
fnc_RTD274 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100010010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(274)
);
fnc_RTD275 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100010011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(275)
);
fnc_RTD276 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100010100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(276)
);
fnc_RTD277 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100010101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(277)
);
fnc_RTD278 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100010110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(278)
);
fnc_RTD279 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100010111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(279)
);
fnc_RTD280 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100011000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(280)
);
fnc_RTD281 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100011001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(281)
);
fnc_RTD282 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100011010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(282)
);
fnc_RTD283 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100011011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(283)
);
fnc_RTD284 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100011100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(284)
);
fnc_RTD285 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100011101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(285)
);
fnc_RTD286 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100011110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(286)
);
fnc_RTD287 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100011111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(287)
);
fnc_RTD288 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100100000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(288)
);
fnc_RTD289 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100100001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(289)
);
fnc_RTD290 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100100010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(290)
);
fnc_RTD291 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100100011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(291)
);
fnc_RTD292 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100100100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(292)
);
fnc_RTD293 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100100101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(293)
);
fnc_RTD294 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100100110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(294)
);
fnc_RTD295 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100100111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(295)
);
fnc_RTD296 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100101000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(296)
);
fnc_RTD297 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100101001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(297)
);
fnc_RTD298 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100101010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(298)
);
fnc_RTD299 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100101011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(299)
);
fnc_RTD300 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100101100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(300)
);
fnc_RTD301 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100101101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(301)
);
fnc_RTD302 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100101110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(302)
);
fnc_RTD303 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100101111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(303)
);
fnc_RTD304 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100110000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(304)
);
fnc_RTD305 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100110001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(305)
);
fnc_RTD306 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100110010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(306)
);
fnc_RTD307 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100110011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(307)
);
fnc_RTD308 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100110100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(308)
);
fnc_RTD309 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100110101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(309)
);
fnc_RTD310 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100110110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(310)
);
fnc_RTD311 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100110111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(311)
);
fnc_RTD312 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100111000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(312)
);
fnc_RTD313 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100111001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(313)
);
fnc_RTD314 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100111010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(314)
);
fnc_RTD315 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100111011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(315)
);
fnc_RTD316 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100111100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(316)
);
fnc_RTD317 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100111101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(317)
);
fnc_RTD318 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100111110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(318)
);
fnc_RTD319 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100111111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(319)
);
fnc_RTD320 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101000000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(320)
);
fnc_RTD321 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101000001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(321)
);
fnc_RTD322 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101000010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(322)
);
fnc_RTD323 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101000011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(323)
);
fnc_RTD324 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101000100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(324)
);
fnc_RTD325 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101000101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(325)
);
fnc_RTD326 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101000110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(326)
);
fnc_RTD327 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101000111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(327)
);
fnc_RTD328 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101001000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(328)
);
fnc_RTD329 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101001001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(329)
);
fnc_RTD330 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101001010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(330)
);
fnc_RTD331 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101001011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(331)
);
fnc_RTD332 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101001100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(332)
);
fnc_RTD333 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101001101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(333)
);
fnc_RTD334 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101001110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(334)
);
fnc_RTD335 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101001111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(335)
);
fnc_RTD336 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101010000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(336)
);
fnc_RTD337 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101010001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(337)
);
fnc_RTD338 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101010010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(338)
);
fnc_RTD339 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101010011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(339)
);
fnc_RTD340 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101010100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(340)
);
fnc_RTD341 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101010101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(341)
);
fnc_RTD342 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101010110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(342)
);
fnc_RTD343 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101010111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(343)
);
fnc_RTD344 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101011000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(344)
);
fnc_RTD345 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101011001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(345)
);
fnc_RTD346 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101011010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(346)
);
fnc_RTD347 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101011011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(347)
);
fnc_RTD348 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101011100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(348)
);
fnc_RTD349 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101011101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(349)
);
fnc_RTD350 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101011110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(350)
);
fnc_RTD351 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101011111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(351)
);
fnc_RTD352 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101100000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(352)
);
fnc_RTD353 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101100001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(353)
);
fnc_RTD354 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101100010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(354)
);
fnc_RTD355 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101100011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(355)
);
fnc_RTD356 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101100100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(356)
);
fnc_RTD357 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101100101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(357)
);
fnc_RTD358 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101100110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(358)
);
fnc_RTD359 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101100111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(359)
);
fnc_RTD360 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101101000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(360)
);
fnc_RTD361 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101101001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(361)
);
fnc_RTD362 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101101010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(362)
);
fnc_RTD363 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101101011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(363)
);
fnc_RTD364 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101101100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(364)
);
fnc_RTD365 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101101101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(365)
);
fnc_RTD366 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101101110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(366)
);
fnc_RTD367 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101101111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(367)
);
fnc_RTD368 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101110000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(368)
);
fnc_RTD369 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101110001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(369)
);
fnc_RTD370 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101110010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(370)
);
fnc_RTD371 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101110011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(371)
);
fnc_RTD372 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101110100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(372)
);
fnc_RTD373 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101110101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(373)
);
fnc_RTD374 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101110110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(374)
);
fnc_RTD375 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101110111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(375)
);
fnc_RTD376 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101111000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(376)
);
fnc_RTD377 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101111001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(377)
);
fnc_RTD378 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101111010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(378)
);
fnc_RTD379 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101111011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(379)
);
fnc_RTD380 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101111100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(380)
);
fnc_RTD381 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101111101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(381)
);
fnc_RTD382 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101111110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(382)
);
fnc_RTD383 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101111111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(383)
);
fnc_RTD384 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110000000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(384)
);
fnc_RTD385 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110000001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(385)
);
fnc_RTD386 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110000010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(386)
);
fnc_RTD387 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110000011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(387)
);
fnc_RTD388 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110000100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(388)
);
fnc_RTD389 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110000101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(389)
);
fnc_RTD390 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110000110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(390)
);
fnc_RTD391 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110000111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(391)
);
fnc_RTD392 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110001000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(392)
);
fnc_RTD393 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110001001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(393)
);
fnc_RTD394 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110001010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(394)
);
fnc_RTD395 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110001011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(395)
);
fnc_RTD396 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110001100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(396)
);
fnc_RTD397 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110001101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(397)
);
fnc_RTD398 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110001110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(398)
);
fnc_RTD399 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110001111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(399)
);
fnc_RTD400 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110010000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(400)
);
fnc_RTD401 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110010001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(401)
);
fnc_RTD402 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110010010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(402)
);
fnc_RTD403 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110010011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(403)
);
fnc_RTD404 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110010100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(404)
);
fnc_RTD405 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110010101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(405)
);
fnc_RTD406 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110010110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(406)
);
fnc_RTD407 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110010111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(407)
);
fnc_RTD408 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110011000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(408)
);
fnc_RTD409 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110011001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(409)
);
fnc_RTD410 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110011010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(410)
);
fnc_RTD411 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110011011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(411)
);
fnc_RTD412 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110011100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(412)
);
fnc_RTD413 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110011101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(413)
);
fnc_RTD414 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110011110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(414)
);
fnc_RTD415 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110011111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(415)
);
fnc_RTD416 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110100000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(416)
);
fnc_RTD417 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110100001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(417)
);
fnc_RTD418 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110100010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(418)
);
fnc_RTD419 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110100011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(419)
);
fnc_RTD420 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110100100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(420)
);
fnc_RTD421 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110100101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(421)
);
fnc_RTD422 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110100110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(422)
);
fnc_RTD423 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110100111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(423)
);
fnc_RTD424 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110101000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(424)
);
fnc_RTD425 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110101001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(425)
);
fnc_RTD426 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110101010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(426)
);
fnc_RTD427 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110101011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(427)
);
fnc_RTD428 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110101100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(428)
);
fnc_RTD429 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110101101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(429)
);
fnc_RTD430 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110101110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(430)
);
fnc_RTD431 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110101111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(431)
);
fnc_RTD432 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110110000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(432)
);
fnc_RTD433 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110110001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(433)
);
fnc_RTD434 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110110010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(434)
);
fnc_RTD435 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110110011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(435)
);
fnc_RTD436 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110110100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(436)
);
fnc_RTD437 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110110101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(437)
);
fnc_RTD438 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110110110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(438)
);
fnc_RTD439 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110110111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(439)
);
fnc_RTD440 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110111000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(440)
);
fnc_RTD441 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110111001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(441)
);
fnc_RTD442 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110111010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(442)
);
fnc_RTD443 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110111011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(443)
);
fnc_RTD444 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110111100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(444)
);
fnc_RTD445 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110111101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(445)
);
fnc_RTD446 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110111110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(446)
);
fnc_RTD447 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110111111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(447)
);
fnc_RTD448 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111000000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(448)
);
fnc_RTD449 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111000001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(449)
);
fnc_RTD450 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111000010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(450)
);
fnc_RTD451 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111000011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(451)
);
fnc_RTD452 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111000100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(452)
);
fnc_RTD453 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111000101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(453)
);
fnc_RTD454 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111000110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(454)
);
fnc_RTD455 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111000111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(455)
);
fnc_RTD456 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111001000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(456)
);
fnc_RTD457 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111001001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(457)
);
fnc_RTD458 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111001010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(458)
);
fnc_RTD459 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111001011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(459)
);
fnc_RTD460 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111001100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(460)
);
fnc_RTD461 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111001101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(461)
);
fnc_RTD462 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111001110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(462)
);
fnc_RTD463 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111001111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(463)
);
fnc_RTD464 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111010000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(464)
);
fnc_RTD465 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111010001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(465)
);
fnc_RTD466 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111010010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(466)
);
fnc_RTD467 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111010011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(467)
);
fnc_RTD468 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111010100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(468)
);
fnc_RTD469 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111010101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(469)
);
fnc_RTD470 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111010110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(470)
);
fnc_RTD471 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111010111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(471)
);
fnc_RTD472 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111011000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(472)
);
fnc_RTD473 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111011001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(473)
);
fnc_RTD474 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111011010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(474)
);
fnc_RTD475 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111011011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(475)
);
fnc_RTD476 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111011100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(476)
);
fnc_RTD477 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111011101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(477)
);
fnc_RTD478 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111011110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(478)
);
fnc_RTD479 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111011111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(479)
);
fnc_RTD480 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111100000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(480)
);
fnc_RTD481 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111100001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(481)
);
fnc_RTD482 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111100010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(482)
);
fnc_RTD483 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111100011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(483)
);
fnc_RTD484 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111100100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(484)
);
fnc_RTD485 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111100101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(485)
);
fnc_RTD486 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111100110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(486)
);
fnc_RTD487 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111100111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(487)
);
fnc_RTD488 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111101000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(488)
);
fnc_RTD489 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111101001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(489)
);
fnc_RTD490 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111101010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(490)
);
fnc_RTD491 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111101011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(491)
);
fnc_RTD492 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111101100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(492)
);
fnc_RTD493 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111101101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(493)
);
fnc_RTD494 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111101110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(494)
);
fnc_RTD495 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111101111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(495)
);
fnc_RTD496 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111110000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(496)
);
fnc_RTD497 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111110001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(497)
);
fnc_RTD498 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111110010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(498)
);
fnc_RTD499 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111110011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(499)
);
fnc_RTD500 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111110100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(500)
);
fnc_RTD501 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111110101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(501)
);
fnc_RTD502 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111110110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(502)
);
fnc_RTD503 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111110111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(503)
);
fnc_RTD504 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111111000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(504)
);
fnc_RTD505 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111111001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(505)
);
fnc_RTD506 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111111010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(506)
);
fnc_RTD507 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111111011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(507)
);
fnc_RTD508 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111111100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(508)
);
fnc_RTD509 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111111101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(509)
);
fnc_RTD510 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111111110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(510)
);
fnc_RTD511 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111111111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(511)
);
fnc_RTD512 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000000000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(512)
);
fnc_RTD513 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000000001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(513)
);
fnc_RTD514 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000000010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(514)
);
fnc_RTD515 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000000011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(515)
);
fnc_RTD516 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000000100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(516)
);
fnc_RTD517 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000000101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(517)
);
fnc_RTD518 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000000110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(518)
);
fnc_RTD519 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000000111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(519)
);
fnc_RTD520 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000001000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(520)
);
fnc_RTD521 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000001001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(521)
);
fnc_RTD522 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000001010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(522)
);
fnc_RTD523 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000001011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(523)
);
fnc_RTD524 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000001100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(524)
);
fnc_RTD525 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000001101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(525)
);
fnc_RTD526 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000001110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(526)
);
fnc_RTD527 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000001111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(527)
);
fnc_RTD528 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000010000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(528)
);
fnc_RTD529 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000010001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(529)
);
fnc_RTD530 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000010010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(530)
);
fnc_RTD531 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000010011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(531)
);
fnc_RTD532 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000010100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(532)
);
fnc_RTD533 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000010101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(533)
);
fnc_RTD534 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000010110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(534)
);
fnc_RTD535 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000010111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(535)
);
fnc_RTD536 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000011000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(536)
);
fnc_RTD537 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000011001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(537)
);
fnc_RTD538 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000011010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(538)
);
fnc_RTD539 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000011011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(539)
);
fnc_RTD540 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000011100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(540)
);
fnc_RTD541 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000011101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(541)
);
fnc_RTD542 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000011110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(542)
);
fnc_RTD543 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000011111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(543)
);
fnc_RTD544 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000100000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(544)
);
fnc_RTD545 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000100001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(545)
);
fnc_RTD546 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000100010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(546)
);
fnc_RTD547 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000100011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(547)
);
fnc_RTD548 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000100100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(548)
);
fnc_RTD549 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000100101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(549)
);
fnc_RTD550 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000100110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(550)
);
fnc_RTD551 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000100111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(551)
);
fnc_RTD552 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000101000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(552)
);
fnc_RTD553 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000101001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(553)
);
fnc_RTD554 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000101010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(554)
);
fnc_RTD555 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000101011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(555)
);
fnc_RTD556 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000101100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(556)
);
fnc_RTD557 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000101101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(557)
);
fnc_RTD558 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000101110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(558)
);
fnc_RTD559 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000101111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(559)
);
fnc_RTD560 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000110000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(560)
);
fnc_RTD561 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000110001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(561)
);
fnc_RTD562 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000110010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(562)
);
fnc_RTD563 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000110011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(563)
);
fnc_RTD564 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000110100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(564)
);
fnc_RTD565 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000110101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(565)
);
fnc_RTD566 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000110110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(566)
);
fnc_RTD567 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000110111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(567)
);
fnc_RTD568 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000111000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(568)
);
fnc_RTD569 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000111001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(569)
);
fnc_RTD570 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000111010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(570)
);
fnc_RTD571 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000111011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(571)
);
fnc_RTD572 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000111100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(572)
);
fnc_RTD573 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000111101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(573)
);
fnc_RTD574 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000111110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(574)
);
fnc_RTD575 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000111111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(575)
);
fnc_RTD576 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001000000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(576)
);
fnc_RTD577 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001000001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(577)
);
fnc_RTD578 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001000010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(578)
);
fnc_RTD579 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001000011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(579)
);
fnc_RTD580 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001000100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(580)
);
fnc_RTD581 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001000101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(581)
);
fnc_RTD582 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001000110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(582)
);
fnc_RTD583 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001000111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(583)
);
fnc_RTD584 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001001000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(584)
);
fnc_RTD585 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001001001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(585)
);
fnc_RTD586 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001001010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(586)
);
fnc_RTD587 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001001011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(587)
);
fnc_RTD588 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001001100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(588)
);
fnc_RTD589 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001001101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(589)
);
fnc_RTD590 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001001110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(590)
);
fnc_RTD591 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001001111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(591)
);
fnc_RTD592 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001010000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(592)
);
fnc_RTD593 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001010001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(593)
);
fnc_RTD594 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001010010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(594)
);
fnc_RTD595 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001010011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(595)
);
fnc_RTD596 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001010100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(596)
);
fnc_RTD597 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001010101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(597)
);
fnc_RTD598 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001010110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(598)
);
fnc_RTD599 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001010111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(599)
);
fnc_RTD600 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001011000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(600)
);
fnc_RTD601 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001011001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(601)
);
fnc_RTD602 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001011010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(602)
);
fnc_RTD603 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001011011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(603)
);
fnc_RTD604 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001011100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(604)
);
fnc_RTD605 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001011101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(605)
);
fnc_RTD606 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001011110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(606)
);
fnc_RTD607 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001011111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(607)
);
fnc_RTD608 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001100000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(608)
);
fnc_RTD609 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001100001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(609)
);
fnc_RTD610 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001100010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(610)
);
fnc_RTD611 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001100011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(611)
);
fnc_RTD612 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001100100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(612)
);
fnc_RTD613 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001100101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(613)
);
fnc_RTD614 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001100110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(614)
);
fnc_RTD615 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001100111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(615)
);
fnc_RTD616 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001101000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(616)
);
fnc_RTD617 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001101001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(617)
);
fnc_RTD618 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001101010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(618)
);
fnc_RTD619 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001101011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(619)
);
fnc_RTD620 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001101100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(620)
);
fnc_RTD621 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001101101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(621)
);
fnc_RTD622 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001101110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(622)
);
fnc_RTD623 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001101111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(623)
);
fnc_RTD624 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001110000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(624)
);
fnc_RTD625 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001110001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(625)
);
fnc_RTD626 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001110010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(626)
);
fnc_RTD627 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001110011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(627)
);
fnc_RTD628 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001110100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(628)
);
fnc_RTD629 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001110101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(629)
);
fnc_RTD630 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001110110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(630)
);
fnc_RTD631 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001110111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(631)
);
fnc_RTD632 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001111000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(632)
);
fnc_RTD633 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001111001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(633)
);
fnc_RTD634 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001111010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(634)
);
fnc_RTD635 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001111011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(635)
);
fnc_RTD636 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001111100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(636)
);
fnc_RTD637 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001111101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(637)
);
fnc_RTD638 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001111110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(638)
);
fnc_RTD639 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001111111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(639)
);
fnc_RTD640 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010000000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(640)
);
fnc_RTD641 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010000001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(641)
);
fnc_RTD642 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010000010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(642)
);
fnc_RTD643 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010000011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(643)
);
fnc_RTD644 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010000100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(644)
);
fnc_RTD645 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010000101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(645)
);
fnc_RTD646 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010000110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(646)
);
fnc_RTD647 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010000111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(647)
);
fnc_RTD648 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010001000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(648)
);
fnc_RTD649 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010001001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(649)
);
fnc_RTD650 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010001010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(650)
);
fnc_RTD651 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010001011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(651)
);
fnc_RTD652 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010001100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(652)
);
fnc_RTD653 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010001101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(653)
);
fnc_RTD654 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010001110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(654)
);
fnc_RTD655 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010001111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(655)
);
fnc_RTD656 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010010000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(656)
);
fnc_RTD657 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010010001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(657)
);
fnc_RTD658 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010010010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(658)
);
fnc_RTD659 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010010011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(659)
);
fnc_RTD660 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010010100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(660)
);
fnc_RTD661 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010010101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(661)
);
fnc_RTD662 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010010110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(662)
);
fnc_RTD663 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010010111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(663)
);
fnc_RTD664 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010011000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(664)
);
fnc_RTD665 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010011001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(665)
);
fnc_RTD666 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010011010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(666)
);
fnc_RTD667 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010011011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(667)
);
fnc_RTD668 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010011100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(668)
);
fnc_RTD669 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010011101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(669)
);
fnc_RTD670 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010011110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(670)
);
fnc_RTD671 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010011111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(671)
);
fnc_RTD672 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010100000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(672)
);
fnc_RTD673 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010100001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(673)
);
fnc_RTD674 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010100010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(674)
);
fnc_RTD675 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010100011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(675)
);
fnc_RTD676 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010100100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(676)
);
fnc_RTD677 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010100101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(677)
);
fnc_RTD678 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010100110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(678)
);
fnc_RTD679 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010100111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(679)
);
fnc_RTD680 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010101000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(680)
);
fnc_RTD681 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010101001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(681)
);
fnc_RTD682 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010101010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(682)
);
fnc_RTD683 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010101011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(683)
);
fnc_RTD684 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010101100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(684)
);
fnc_RTD685 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010101101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(685)
);
fnc_RTD686 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010101110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(686)
);
fnc_RTD687 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010101111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(687)
);
fnc_RTD688 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010110000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(688)
);
fnc_RTD689 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010110001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(689)
);
fnc_RTD690 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010110010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(690)
);
fnc_RTD691 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010110011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(691)
);
fnc_RTD692 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010110100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(692)
);
fnc_RTD693 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010110101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(693)
);
fnc_RTD694 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010110110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(694)
);
fnc_RTD695 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010110111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(695)
);
fnc_RTD696 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010111000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(696)
);
fnc_RTD697 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010111001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(697)
);
fnc_RTD698 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010111010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(698)
);
fnc_RTD699 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010111011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(699)
);
fnc_RTD700 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010111100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(700)
);
fnc_RTD701 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010111101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(701)
);
fnc_RTD702 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010111110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(702)
);
fnc_RTD703 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010111111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(703)
);
fnc_RTD704 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011000000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(704)
);
fnc_RTD705 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011000001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(705)
);
fnc_RTD706 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011000010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(706)
);
fnc_RTD707 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011000011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(707)
);
fnc_RTD708 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011000100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(708)
);
fnc_RTD709 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011000101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(709)
);
fnc_RTD710 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011000110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(710)
);
fnc_RTD711 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011000111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(711)
);
fnc_RTD712 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011001000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(712)
);
fnc_RTD713 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011001001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(713)
);
fnc_RTD714 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011001010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(714)
);
fnc_RTD715 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011001011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(715)
);
fnc_RTD716 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011001100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(716)
);
fnc_RTD717 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011001101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(717)
);
fnc_RTD718 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011001110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(718)
);
fnc_RTD719 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011001111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(719)
);
fnc_RTD720 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011010000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(720)
);
fnc_RTD721 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011010001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(721)
);
fnc_RTD722 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011010010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(722)
);
fnc_RTD723 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011010011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(723)
);
fnc_RTD724 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011010100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(724)
);
fnc_RTD725 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011010101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(725)
);
fnc_RTD726 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011010110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(726)
);
fnc_RTD727 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011010111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(727)
);
fnc_RTD728 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011011000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(728)
);
fnc_RTD729 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011011001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(729)
);
fnc_RTD730 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011011010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(730)
);
fnc_RTD731 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011011011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(731)
);
fnc_RTD732 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011011100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(732)
);
fnc_RTD733 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011011101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(733)
);
fnc_RTD734 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011011110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(734)
);
fnc_RTD735 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011011111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(735)
);
fnc_RTD736 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011100000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(736)
);
fnc_RTD737 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011100001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(737)
);
fnc_RTD738 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011100010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(738)
);
fnc_RTD739 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011100011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(739)
);
fnc_RTD740 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011100100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(740)
);
fnc_RTD741 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011100101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(741)
);
fnc_RTD742 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011100110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(742)
);
fnc_RTD743 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011100111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(743)
);
fnc_RTD744 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011101000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(744)
);
fnc_RTD745 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011101001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(745)
);
fnc_RTD746 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011101010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(746)
);
fnc_RTD747 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011101011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(747)
);
fnc_RTD748 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011101100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(748)
);
fnc_RTD749 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011101101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(749)
);
fnc_RTD750 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011101110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(750)
);
fnc_RTD751 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011101111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(751)
);
fnc_RTD752 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011110000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(752)
);
fnc_RTD753 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011110001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(753)
);
fnc_RTD754 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011110010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(754)
);
fnc_RTD755 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011110011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(755)
);
fnc_RTD756 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011110100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(756)
);
fnc_RTD757 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011110101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(757)
);
fnc_RTD758 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011110110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(758)
);
fnc_RTD759 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011110111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(759)
);
fnc_RTD760 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011111000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(760)
);
fnc_RTD761 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011111001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(761)
);
fnc_RTD762 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011111010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(762)
);
fnc_RTD763 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011111011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(763)
);
fnc_RTD764 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011111100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(764)
);
fnc_RTD765 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011111101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(765)
);
fnc_RTD766 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011111110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(766)
);
fnc_RTD767 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011111111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(767)
);
fnc_RTD768 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100000000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(768)
);
fnc_RTD769 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100000001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(769)
);
fnc_RTD770 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100000010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(770)
);
fnc_RTD771 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100000011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(771)
);
fnc_RTD772 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100000100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(772)
);
fnc_RTD773 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100000101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(773)
);
fnc_RTD774 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100000110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(774)
);
fnc_RTD775 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100000111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(775)
);
fnc_RTD776 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100001000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(776)
);
fnc_RTD777 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100001001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(777)
);
fnc_RTD778 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100001010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(778)
);
fnc_RTD779 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100001011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(779)
);
fnc_RTD780 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100001100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(780)
);
fnc_RTD781 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100001101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(781)
);
fnc_RTD782 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100001110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(782)
);
fnc_RTD783 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100001111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(783)
);
fnc_RTD784 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100010000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(784)
);
fnc_RTD785 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100010001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(785)
);
fnc_RTD786 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100010010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(786)
);
fnc_RTD787 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100010011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(787)
);
fnc_RTD788 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100010100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(788)
);
fnc_RTD789 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100010101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(789)
);
fnc_RTD790 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100010110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(790)
);
fnc_RTD791 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100010111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(791)
);
fnc_RTD792 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100011000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(792)
);
fnc_RTD793 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100011001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(793)
);
fnc_RTD794 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100011010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(794)
);
fnc_RTD795 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100011011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(795)
);
fnc_RTD796 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100011100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(796)
);
fnc_RTD797 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100011101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(797)
);
fnc_RTD798 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100011110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(798)
);
fnc_RTD799 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100011111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(799)
);
fnc_RTD800 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100100000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(800)
);
fnc_RTD801 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100100001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(801)
);
fnc_RTD802 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100100010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(802)
);
fnc_RTD803 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100100011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(803)
);
fnc_RTD804 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100100100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(804)
);
fnc_RTD805 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100100101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(805)
);
fnc_RTD806 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100100110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(806)
);
fnc_RTD807 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100100111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(807)
);
fnc_RTD808 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100101000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(808)
);
fnc_RTD809 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100101001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(809)
);
fnc_RTD810 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100101010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(810)
);
fnc_RTD811 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100101011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(811)
);
fnc_RTD812 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100101100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(812)
);
fnc_RTD813 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100101101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(813)
);
fnc_RTD814 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100101110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(814)
);
fnc_RTD815 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100101111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(815)
);
fnc_RTD816 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100110000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(816)
);
fnc_RTD817 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100110001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(817)
);
fnc_RTD818 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100110010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(818)
);
fnc_RTD819 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100110011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(819)
);
fnc_RTD820 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100110100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(820)
);
fnc_RTD821 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100110101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(821)
);
fnc_RTD822 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100110110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(822)
);
fnc_RTD823 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100110111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(823)
);
fnc_RTD824 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100111000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(824)
);
fnc_RTD825 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100111001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(825)
);
fnc_RTD826 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100111010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(826)
);
fnc_RTD827 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100111011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(827)
);
fnc_RTD828 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100111100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(828)
);
fnc_RTD829 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100111101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(829)
);
fnc_RTD830 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100111110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(830)
);
fnc_RTD831 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100111111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(831)
);
fnc_RTD832 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101000000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(832)
);
fnc_RTD833 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101000001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(833)
);
fnc_RTD834 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101000010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(834)
);
fnc_RTD835 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101000011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(835)
);
fnc_RTD836 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101000100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(836)
);
fnc_RTD837 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101000101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(837)
);
fnc_RTD838 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101000110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(838)
);
fnc_RTD839 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101000111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(839)
);
fnc_RTD840 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101001000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(840)
);
fnc_RTD841 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101001001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(841)
);
fnc_RTD842 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101001010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(842)
);
fnc_RTD843 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101001011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(843)
);
fnc_RTD844 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101001100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(844)
);
fnc_RTD845 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101001101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(845)
);
fnc_RTD846 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101001110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(846)
);
fnc_RTD847 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101001111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(847)
);
fnc_RTD848 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101010000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(848)
);
fnc_RTD849 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101010001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(849)
);
fnc_RTD850 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101010010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(850)
);
fnc_RTD851 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101010011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(851)
);
fnc_RTD852 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101010100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(852)
);
fnc_RTD853 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101010101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(853)
);
fnc_RTD854 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101010110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(854)
);
fnc_RTD855 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101010111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(855)
);
fnc_RTD856 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101011000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(856)
);
fnc_RTD857 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101011001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(857)
);
fnc_RTD858 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101011010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(858)
);
fnc_RTD859 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101011011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(859)
);
fnc_RTD860 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101011100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(860)
);
fnc_RTD861 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101011101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(861)
);
fnc_RTD862 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101011110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(862)
);
fnc_RTD863 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101011111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(863)
);
fnc_RTD864 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101100000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(864)
);
fnc_RTD865 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101100001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(865)
);
fnc_RTD866 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101100010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(866)
);
fnc_RTD867 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101100011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(867)
);
fnc_RTD868 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101100100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(868)
);
fnc_RTD869 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101100101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(869)
);
fnc_RTD870 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101100110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(870)
);
fnc_RTD871 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101100111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(871)
);
fnc_RTD872 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101101000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(872)
);
fnc_RTD873 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101101001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(873)
);
fnc_RTD874 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101101010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(874)
);
fnc_RTD875 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101101011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(875)
);
fnc_RTD876 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101101100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(876)
);
fnc_RTD877 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101101101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(877)
);
fnc_RTD878 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101101110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(878)
);
fnc_RTD879 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101101111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(879)
);
fnc_RTD880 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101110000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(880)
);
fnc_RTD881 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101110001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(881)
);
fnc_RTD882 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101110010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(882)
);
fnc_RTD883 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101110011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(883)
);
fnc_RTD884 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101110100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(884)
);
fnc_RTD885 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101110101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(885)
);
fnc_RTD886 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101110110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(886)
);
fnc_RTD887 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101110111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(887)
);
fnc_RTD888 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101111000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(888)
);
fnc_RTD889 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101111001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(889)
);
fnc_RTD890 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101111010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(890)
);
fnc_RTD891 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101111011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(891)
);
fnc_RTD892 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101111100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(892)
);
fnc_RTD893 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101111101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(893)
);
fnc_RTD894 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101111110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(894)
);
fnc_RTD895 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101111111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(895)
);
fnc_RTD896 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110000000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(896)
);
fnc_RTD897 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110000001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(897)
);
fnc_RTD898 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110000010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(898)
);
fnc_RTD899 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110000011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(899)
);
fnc_RTD900 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110000100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(900)
);
fnc_RTD901 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110000101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(901)
);
fnc_RTD902 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110000110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(902)
);
fnc_RTD903 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110000111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(903)
);
fnc_RTD904 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110001000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(904)
);
fnc_RTD905 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110001001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(905)
);
fnc_RTD906 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110001010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(906)
);
fnc_RTD907 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110001011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(907)
);
fnc_RTD908 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110001100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(908)
);
fnc_RTD909 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110001101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(909)
);
fnc_RTD910 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110001110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(910)
);
fnc_RTD911 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110001111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(911)
);
fnc_RTD912 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110010000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(912)
);
fnc_RTD913 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110010001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(913)
);
fnc_RTD914 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110010010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(914)
);
fnc_RTD915 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110010011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(915)
);
fnc_RTD916 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110010100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(916)
);
fnc_RTD917 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110010101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(917)
);
fnc_RTD918 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110010110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(918)
);
fnc_RTD919 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110010111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(919)
);
fnc_RTD920 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110011000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(920)
);
fnc_RTD921 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110011001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(921)
);
fnc_RTD922 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110011010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(922)
);
fnc_RTD923 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110011011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(923)
);
fnc_RTD924 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110011100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(924)
);
fnc_RTD925 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110011101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(925)
);
fnc_RTD926 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110011110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(926)
);
fnc_RTD927 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110011111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(927)
);
fnc_RTD928 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110100000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(928)
);
fnc_RTD929 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110100001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(929)
);
fnc_RTD930 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110100010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(930)
);
fnc_RTD931 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110100011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(931)
);
fnc_RTD932 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110100100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(932)
);
fnc_RTD933 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110100101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(933)
);
fnc_RTD934 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110100110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(934)
);
fnc_RTD935 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110100111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(935)
);
fnc_RTD936 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110101000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(936)
);
fnc_RTD937 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110101001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(937)
);
fnc_RTD938 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110101010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(938)
);
fnc_RTD939 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110101011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(939)
);
fnc_RTD940 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110101100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(940)
);
fnc_RTD941 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110101101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(941)
);
fnc_RTD942 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110101110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(942)
);
fnc_RTD943 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110101111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(943)
);
fnc_RTD944 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110110000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(944)
);
fnc_RTD945 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110110001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(945)
);
fnc_RTD946 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110110010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(946)
);
fnc_RTD947 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110110011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(947)
);
fnc_RTD948 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110110100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(948)
);
fnc_RTD949 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110110101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(949)
);
fnc_RTD950 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110110110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(950)
);
fnc_RTD951 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110110111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(951)
);
fnc_RTD952 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110111000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(952)
);
fnc_RTD953 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110111001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(953)
);
fnc_RTD954 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110111010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(954)
);
fnc_RTD955 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110111011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(955)
);
fnc_RTD956 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110111100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(956)
);
fnc_RTD957 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110111101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(957)
);
fnc_RTD958 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110111110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(958)
);
fnc_RTD959 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110111111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(959)
);
fnc_RTD960 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111000000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(960)
);
fnc_RTD961 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111000001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(961)
);
fnc_RTD962 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111000010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(962)
);
fnc_RTD963 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111000011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(963)
);
fnc_RTD964 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111000100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(964)
);
fnc_RTD965 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111000101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(965)
);
fnc_RTD966 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111000110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(966)
);
fnc_RTD967 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111000111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(967)
);
fnc_RTD968 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111001000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(968)
);
fnc_RTD969 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111001001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(969)
);
fnc_RTD970 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111001010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(970)
);
fnc_RTD971 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111001011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(971)
);
fnc_RTD972 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111001100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(972)
);
fnc_RTD973 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111001101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(973)
);
fnc_RTD974 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111001110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(974)
);
fnc_RTD975 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111001111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(975)
);
fnc_RTD976 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111010000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(976)
);
fnc_RTD977 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111010001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(977)
);
fnc_RTD978 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111010010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(978)
);
fnc_RTD979 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111010011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(979)
);
fnc_RTD980 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111010100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(980)
);
fnc_RTD981 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111010101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(981)
);
fnc_RTD982 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111010110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(982)
);
fnc_RTD983 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111010111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(983)
);
fnc_RTD984 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111011000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(984)
);
fnc_RTD985 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111011001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(985)
);
fnc_RTD986 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111011010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(986)
);
fnc_RTD987 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111011011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(987)
);
fnc_RTD988 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111011100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(988)
);
fnc_RTD989 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111011101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(989)
);
fnc_RTD990 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111011110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(990)
);
fnc_RTD991 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111011111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(991)
);
fnc_RTD992 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111100000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(992)
);
fnc_RTD993 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111100001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(993)
);
fnc_RTD994 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111100010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(994)
);
fnc_RTD995 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111100011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(995)
);
fnc_RTD996 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111100100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(996)
);
fnc_RTD997 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111100101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(997)
);
fnc_RTD998 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111100110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(998)
);
fnc_RTD999 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111100111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(999)
);
fnc_RTD1000 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111101000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1000)
);
fnc_RTD1001 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111101001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1001)
);
fnc_RTD1002 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111101010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1002)
);
fnc_RTD1003 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111101011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1003)
);
fnc_RTD1004 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111101100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1004)
);
fnc_RTD1005 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111101101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1005)
);
fnc_RTD1006 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111101110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1006)
);
fnc_RTD1007 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111101111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1007)
);
fnc_RTD1008 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111110000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1008)
);
fnc_RTD1009 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111110001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1009)
);
fnc_RTD1010 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111110010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1010)
);
fnc_RTD1011 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111110011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1011)
);
fnc_RTD1012 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111110100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1012)
);
fnc_RTD1013 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111110101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1013)
);
fnc_RTD1014 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111110110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1014)
);
fnc_RTD1015 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111110111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1015)
);
fnc_RTD1016 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111111000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1016)
);
fnc_RTD1017 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111111001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1017)
);
fnc_RTD1018 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111111010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1018)
);
fnc_RTD1019 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111111011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1019)
);
fnc_RTD1020 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111111100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1020)
);
fnc_RTD1021 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111111101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1021)
);
fnc_RTD1022 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111111110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1022)
);
fnc_RTD1023 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111111111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1023)
);
fnc_RTD1024 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000000000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1024)
);
fnc_RTD1025 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000000001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1025)
);
fnc_RTD1026 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000000010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1026)
);
fnc_RTD1027 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000000011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1027)
);
fnc_RTD1028 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000000100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1028)
);
fnc_RTD1029 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000000101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1029)
);
fnc_RTD1030 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000000110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1030)
);
fnc_RTD1031 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000000111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1031)
);
fnc_RTD1032 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000001000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1032)
);
fnc_RTD1033 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000001001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1033)
);
fnc_RTD1034 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000001010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1034)
);
fnc_RTD1035 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000001011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1035)
);
fnc_RTD1036 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000001100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1036)
);
fnc_RTD1037 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000001101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1037)
);
fnc_RTD1038 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000001110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1038)
);
fnc_RTD1039 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000001111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1039)
);
fnc_RTD1040 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000010000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1040)
);
fnc_RTD1041 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000010001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1041)
);
fnc_RTD1042 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000010010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1042)
);
fnc_RTD1043 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000010011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1043)
);
fnc_RTD1044 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000010100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1044)
);
fnc_RTD1045 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000010101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1045)
);
fnc_RTD1046 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000010110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1046)
);
fnc_RTD1047 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000010111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1047)
);
fnc_RTD1048 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000011000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1048)
);
fnc_RTD1049 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000011001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1049)
);
fnc_RTD1050 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000011010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1050)
);
fnc_RTD1051 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000011011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1051)
);
fnc_RTD1052 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000011100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1052)
);
fnc_RTD1053 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000011101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1053)
);
fnc_RTD1054 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000011110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1054)
);
fnc_RTD1055 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000011111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1055)
);
fnc_RTD1056 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000100000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1056)
);
fnc_RTD1057 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000100001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1057)
);
fnc_RTD1058 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000100010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1058)
);
fnc_RTD1059 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000100011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1059)
);
fnc_RTD1060 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000100100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1060)
);
fnc_RTD1061 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000100101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1061)
);
fnc_RTD1062 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000100110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1062)
);
fnc_RTD1063 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000100111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1063)
);
fnc_RTD1064 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000101000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1064)
);
fnc_RTD1065 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000101001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1065)
);
fnc_RTD1066 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000101010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1066)
);
fnc_RTD1067 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000101011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1067)
);
fnc_RTD1068 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000101100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1068)
);
fnc_RTD1069 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000101101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1069)
);
fnc_RTD1070 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000101110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1070)
);
fnc_RTD1071 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000101111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1071)
);
fnc_RTD1072 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000110000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1072)
);
fnc_RTD1073 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000110001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1073)
);
fnc_RTD1074 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000110010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1074)
);
fnc_RTD1075 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000110011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1075)
);
fnc_RTD1076 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000110100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1076)
);
fnc_RTD1077 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000110101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1077)
);
fnc_RTD1078 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000110110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1078)
);
fnc_RTD1079 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000110111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1079)
);
fnc_RTD1080 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000111000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1080)
);
fnc_RTD1081 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000111001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1081)
);
fnc_RTD1082 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000111010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1082)
);
fnc_RTD1083 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000111011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1083)
);
fnc_RTD1084 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000111100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1084)
);
fnc_RTD1085 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000111101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1085)
);
fnc_RTD1086 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000111110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1086)
);
fnc_RTD1087 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000111111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1087)
);
fnc_RTD1088 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001000000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1088)
);
fnc_RTD1089 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001000001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1089)
);
fnc_RTD1090 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001000010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1090)
);
fnc_RTD1091 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001000011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1091)
);
fnc_RTD1092 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001000100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1092)
);
fnc_RTD1093 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001000101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1093)
);
fnc_RTD1094 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001000110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1094)
);
fnc_RTD1095 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001000111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1095)
);
fnc_RTD1096 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001001000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1096)
);
fnc_RTD1097 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001001001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1097)
);
fnc_RTD1098 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001001010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1098)
);
fnc_RTD1099 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001001011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1099)
);
fnc_RTD1100 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001001100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1100)
);
fnc_RTD1101 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001001101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1101)
);
fnc_RTD1102 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001001110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1102)
);
fnc_RTD1103 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001001111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1103)
);
fnc_RTD1104 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001010000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1104)
);
fnc_RTD1105 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001010001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1105)
);
fnc_RTD1106 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001010010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1106)
);
fnc_RTD1107 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001010011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1107)
);
fnc_RTD1108 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001010100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1108)
);
fnc_RTD1109 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001010101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1109)
);
fnc_RTD1110 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001010110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1110)
);
fnc_RTD1111 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001010111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1111)
);
fnc_RTD1112 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001011000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1112)
);
fnc_RTD1113 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001011001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1113)
);
fnc_RTD1114 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001011010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1114)
);
fnc_RTD1115 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001011011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1115)
);
fnc_RTD1116 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001011100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1116)
);
fnc_RTD1117 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001011101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1117)
);
fnc_RTD1118 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001011110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1118)
);
fnc_RTD1119 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001011111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1119)
);
fnc_RTD1120 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001100000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1120)
);
fnc_RTD1121 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001100001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1121)
);
fnc_RTD1122 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001100010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1122)
);
fnc_RTD1123 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001100011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1123)
);
fnc_RTD1124 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001100100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1124)
);
fnc_RTD1125 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001100101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1125)
);
fnc_RTD1126 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001100110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1126)
);
fnc_RTD1127 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001100111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1127)
);
fnc_RTD1128 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001101000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1128)
);
fnc_RTD1129 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001101001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1129)
);
fnc_RTD1130 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001101010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1130)
);
fnc_RTD1131 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001101011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1131)
);
fnc_RTD1132 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001101100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1132)
);
fnc_RTD1133 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001101101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1133)
);
fnc_RTD1134 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001101110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1134)
);
fnc_RTD1135 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001101111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1135)
);
fnc_RTD1136 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001110000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1136)
);
fnc_RTD1137 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001110001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1137)
);
fnc_RTD1138 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001110010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1138)
);
fnc_RTD1139 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001110011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1139)
);
fnc_RTD1140 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001110100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1140)
);
fnc_RTD1141 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001110101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1141)
);
fnc_RTD1142 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001110110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1142)
);
fnc_RTD1143 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001110111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1143)
);
fnc_RTD1144 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001111000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1144)
);
fnc_RTD1145 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001111001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1145)
);
fnc_RTD1146 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001111010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1146)
);
fnc_RTD1147 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001111011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1147)
);
fnc_RTD1148 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001111100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1148)
);
fnc_RTD1149 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001111101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1149)
);
fnc_RTD1150 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001111110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1150)
);
fnc_RTD1151 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001111111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1151)
);
fnc_RTD1152 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010000000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1152)
);
fnc_RTD1153 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010000001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1153)
);
fnc_RTD1154 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010000010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1154)
);
fnc_RTD1155 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010000011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1155)
);
fnc_RTD1156 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010000100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1156)
);
fnc_RTD1157 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010000101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1157)
);
fnc_RTD1158 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010000110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1158)
);
fnc_RTD1159 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010000111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1159)
);
fnc_RTD1160 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010001000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1160)
);
fnc_RTD1161 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010001001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1161)
);
fnc_RTD1162 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010001010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1162)
);
fnc_RTD1163 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010001011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1163)
);
fnc_RTD1164 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010001100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1164)
);
fnc_RTD1165 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010001101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1165)
);
fnc_RTD1166 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010001110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1166)
);
fnc_RTD1167 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010001111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1167)
);
fnc_RTD1168 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010010000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1168)
);
fnc_RTD1169 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010010001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1169)
);
fnc_RTD1170 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010010010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1170)
);
fnc_RTD1171 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010010011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1171)
);
fnc_RTD1172 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010010100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1172)
);
fnc_RTD1173 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010010101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1173)
);
fnc_RTD1174 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010010110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1174)
);
fnc_RTD1175 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010010111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1175)
);
fnc_RTD1176 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010011000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1176)
);
fnc_RTD1177 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010011001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1177)
);
fnc_RTD1178 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010011010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1178)
);
fnc_RTD1179 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010011011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1179)
);
fnc_RTD1180 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010011100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1180)
);
fnc_RTD1181 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010011101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1181)
);
fnc_RTD1182 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010011110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1182)
);
fnc_RTD1183 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010011111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1183)
);
fnc_RTD1184 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010100000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1184)
);
fnc_RTD1185 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010100001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1185)
);
fnc_RTD1186 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010100010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1186)
);
fnc_RTD1187 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010100011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1187)
);
fnc_RTD1188 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010100100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1188)
);
fnc_RTD1189 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010100101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1189)
);
fnc_RTD1190 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010100110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1190)
);
fnc_RTD1191 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010100111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1191)
);
fnc_RTD1192 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010101000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1192)
);
fnc_RTD1193 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010101001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1193)
);
fnc_RTD1194 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010101010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1194)
);
fnc_RTD1195 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010101011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1195)
);
fnc_RTD1196 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010101100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1196)
);
fnc_RTD1197 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010101101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1197)
);
fnc_RTD1198 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010101110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1198)
);
fnc_RTD1199 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010101111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1199)
);
fnc_RTD1200 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010110000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1200)
);
fnc_RTD1201 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010110001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1201)
);
fnc_RTD1202 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010110010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1202)
);
fnc_RTD1203 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010110011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1203)
);
fnc_RTD1204 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010110100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1204)
);
fnc_RTD1205 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010110101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1205)
);
fnc_RTD1206 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010110110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1206)
);
fnc_RTD1207 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010110111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1207)
);
fnc_RTD1208 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010111000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1208)
);
fnc_RTD1209 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010111001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1209)
);
fnc_RTD1210 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010111010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1210)
);
fnc_RTD1211 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010111011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1211)
);
fnc_RTD1212 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010111100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1212)
);
fnc_RTD1213 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010111101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1213)
);
fnc_RTD1214 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010111110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1214)
);
fnc_RTD1215 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010111111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1215)
);
fnc_RTD1216 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010011000000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1216)
);
fnc_RTD1217 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010011000001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1217)
);
fnc_RTD1218 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010011000010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1218)
);
fnc_RTD1219 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010011000011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1219)
);
fnc_RTD1220 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010011000100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1220)
);
fnc_RTD1221 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010011000101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1221)
);
fnc_RTD1222 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010011000110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1222)
);
fnc_RTD1223 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010011000111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1223)
);
fnc_RTD1224 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010011001000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1224)
);
fnc_RTD1225 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010011001001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1225)
);
fnc_RTD1226 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010011001010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1226)
);
fnc_RTD1227 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010011001011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1227)
);
fnc_RTD1228 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010011001100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1228)
);
fnc_RTD1229 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010011001101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1229)
);
fnc_RTD1230 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010011001110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1230)
);
fnc_RTD1231 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010011001111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1231)
);
fnc_RTD1232 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010011010000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1232)
);
fnc_RTD1233 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010011010001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1233)
);
fnc_RTD1234 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010011010010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1234)
);
fnc_RTD1235 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010011010011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1235)
);
fnc_RTD1236 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010011010100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1236)
);
fnc_RTD1237 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010011010101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1237)
);
fnc_RTD1238 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010011010110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1238)
);
fnc_RTD1239 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010011010111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1239)
);
fnc_RTD1240 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010011011000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1240)
);
fnc_RTD1241 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010011011001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1241)
);
fnc_RTD1242 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010011011010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1242)
);
fnc_RTD1243 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010011011011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1243)
);
fnc_RTD1244 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010011011100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1244)
);
fnc_RTD1245 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010011011101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1245)
);
fnc_RTD1246 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010011011110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1246)
);
fnc_RTD1247 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010011011111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1247)
);
fnc_RTD1248 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010011100000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1248)
);
fnc_RTD1249 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010011100001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1249)
);
fnc_RTD1250 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010011100010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1250)
);
fnc_RTD1251 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010011100011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1251)
);
fnc_RTD1252 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010011100100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1252)
);
fnc_RTD1253 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010011100101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1253)
);
fnc_RTD1254 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010011100110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1254)
);
fnc_RTD1255 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010011100111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1255)
);
fnc_RTD1256 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010011101000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1256)
);
fnc_RTD1257 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010011101001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1257)
);
fnc_RTD1258 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010011101010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1258)
);
fnc_RTD1259 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010011101011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1259)
);
fnc_RTD1260 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010011101100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1260)
);
fnc_RTD1261 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010011101101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1261)
);
fnc_RTD1262 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010011101110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1262)
);
fnc_RTD1263 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010011101111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1263)
);
fnc_RTD1264 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010011110000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1264)
);
fnc_RTD1265 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010011110001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1265)
);
fnc_RTD1266 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010011110010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1266)
);
fnc_RTD1267 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010011110011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1267)
);
fnc_RTD1268 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010011110100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1268)
);
fnc_RTD1269 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010011110101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1269)
);
fnc_RTD1270 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010011110110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1270)
);
fnc_RTD1271 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010011110111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1271)
);
fnc_RTD1272 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010011111000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1272)
);
fnc_RTD1273 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010011111001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1273)
);
fnc_RTD1274 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010011111010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1274)
);
fnc_RTD1275 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010011111011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1275)
);
fnc_RTD1276 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010011111100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1276)
);
fnc_RTD1277 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010011111101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1277)
);
fnc_RTD1278 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010011111110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1278)
);
fnc_RTD1279 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010011111111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1279)
);
fnc_RTD1280 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010100000000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1280)
);
fnc_RTD1281 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010100000001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1281)
);
fnc_RTD1282 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010100000010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1282)
);
fnc_RTD1283 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010100000011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1283)
);
fnc_RTD1284 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010100000100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1284)
);
fnc_RTD1285 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010100000101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1285)
);
fnc_RTD1286 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010100000110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1286)
);
fnc_RTD1287 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010100000111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1287)
);
fnc_RTD1288 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010100001000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1288)
);
fnc_RTD1289 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010100001001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1289)
);
fnc_RTD1290 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010100001010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1290)
);
fnc_RTD1291 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010100001011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1291)
);
fnc_RTD1292 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010100001100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1292)
);
fnc_RTD1293 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010100001101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1293)
);
fnc_RTD1294 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010100001110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1294)
);
fnc_RTD1295 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010100001111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1295)
);
fnc_RTD1296 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010100010000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1296)
);
fnc_RTD1297 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010100010001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1297)
);
fnc_RTD1298 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010100010010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1298)
);
fnc_RTD1299 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010100010011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1299)
);
fnc_RTD1300 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010100010100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1300)
);
fnc_RTD1301 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010100010101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1301)
);
fnc_RTD1302 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010100010110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1302)
);
fnc_RTD1303 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010100010111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1303)
);
fnc_RTD1304 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010100011000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1304)
);
fnc_RTD1305 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010100011001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1305)
);
fnc_RTD1306 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010100011010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1306)
);
fnc_RTD1307 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010100011011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1307)
);
fnc_RTD1308 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010100011100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1308)
);
fnc_RTD1309 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010100011101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1309)
);
fnc_RTD1310 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010100011110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1310)
);
fnc_RTD1311 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010100011111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1311)
);
fnc_RTD1312 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010100100000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1312)
);
fnc_RTD1313 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010100100001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1313)
);
fnc_RTD1314 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010100100010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1314)
);
fnc_RTD1315 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010100100011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1315)
);
fnc_RTD1316 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010100100100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1316)
);
fnc_RTD1317 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010100100101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1317)
);
fnc_RTD1318 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010100100110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1318)
);
fnc_RTD1319 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010100100111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1319)
);
fnc_RTD1320 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010100101000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1320)
);
fnc_RTD1321 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010100101001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1321)
);
fnc_RTD1322 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010100101010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1322)
);
fnc_RTD1323 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010100101011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1323)
);
fnc_RTD1324 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010100101100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1324)
);
fnc_RTD1325 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010100101101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1325)
);
fnc_RTD1326 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010100101110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1326)
);
fnc_RTD1327 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010100101111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1327)
);
fnc_RTD1328 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010100110000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1328)
);
fnc_RTD1329 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010100110001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1329)
);
fnc_RTD1330 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010100110010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1330)
);
fnc_RTD1331 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010100110011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1331)
);
fnc_RTD1332 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010100110100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1332)
);
fnc_RTD1333 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010100110101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1333)
);
fnc_RTD1334 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010100110110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1334)
);
fnc_RTD1335 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010100110111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1335)
);
fnc_RTD1336 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010100111000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1336)
);
fnc_RTD1337 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010100111001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1337)
);
fnc_RTD1338 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010100111010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1338)
);
fnc_RTD1339 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010100111011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1339)
);
fnc_RTD1340 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010100111100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1340)
);
fnc_RTD1341 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010100111101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1341)
);
fnc_RTD1342 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010100111110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1342)
);
fnc_RTD1343 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010100111111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1343)
);
fnc_RTD1344 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010101000000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1344)
);
fnc_RTD1345 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010101000001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1345)
);
fnc_RTD1346 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010101000010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1346)
);
fnc_RTD1347 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010101000011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1347)
);
fnc_RTD1348 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010101000100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1348)
);
fnc_RTD1349 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010101000101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1349)
);
fnc_RTD1350 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010101000110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1350)
);
fnc_RTD1351 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010101000111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1351)
);
fnc_RTD1352 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010101001000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1352)
);
fnc_RTD1353 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010101001001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1353)
);
fnc_RTD1354 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010101001010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1354)
);
fnc_RTD1355 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010101001011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1355)
);
fnc_RTD1356 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010101001100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1356)
);
fnc_RTD1357 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010101001101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1357)
);
fnc_RTD1358 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010101001110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1358)
);
fnc_RTD1359 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010101001111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1359)
);
fnc_RTD1360 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010101010000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1360)
);
fnc_RTD1361 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010101010001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1361)
);
fnc_RTD1362 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010101010010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1362)
);
fnc_RTD1363 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010101010011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1363)
);
fnc_RTD1364 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010101010100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1364)
);
fnc_RTD1365 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010101010101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1365)
);
fnc_RTD1366 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010101010110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1366)
);
fnc_RTD1367 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010101010111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1367)
);
fnc_RTD1368 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010101011000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1368)
);
fnc_RTD1369 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010101011001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1369)
);
fnc_RTD1370 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010101011010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1370)
);
fnc_RTD1371 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010101011011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1371)
);
fnc_RTD1372 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010101011100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1372)
);
fnc_RTD1373 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010101011101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1373)
);
fnc_RTD1374 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010101011110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1374)
);
fnc_RTD1375 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010101011111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1375)
);
fnc_RTD1376 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010101100000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1376)
);
fnc_RTD1377 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010101100001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1377)
);
fnc_RTD1378 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010101100010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1378)
);
fnc_RTD1379 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010101100011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1379)
);
fnc_RTD1380 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010101100100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1380)
);
fnc_RTD1381 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010101100101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1381)
);
fnc_RTD1382 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010101100110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1382)
);
fnc_RTD1383 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010101100111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1383)
);
fnc_RTD1384 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010101101000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1384)
);
fnc_RTD1385 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010101101001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1385)
);
fnc_RTD1386 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010101101010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1386)
);
fnc_RTD1387 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010101101011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1387)
);
fnc_RTD1388 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010101101100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1388)
);
fnc_RTD1389 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010101101101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1389)
);
fnc_RTD1390 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010101101110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1390)
);
fnc_RTD1391 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010101101111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1391)
);
fnc_RTD1392 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010101110000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1392)
);
fnc_RTD1393 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010101110001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1393)
);
fnc_RTD1394 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010101110010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1394)
);
fnc_RTD1395 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010101110011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1395)
);
fnc_RTD1396 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010101110100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1396)
);
fnc_RTD1397 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010101110101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1397)
);
fnc_RTD1398 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010101110110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1398)
);
fnc_RTD1399 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010101110111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1399)
);
fnc_RTD1400 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010101111000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1400)
);
fnc_RTD1401 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010101111001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1401)
);
fnc_RTD1402 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010101111010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1402)
);
fnc_RTD1403 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010101111011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1403)
);
fnc_RTD1404 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010101111100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1404)
);
fnc_RTD1405 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010101111101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1405)
);
fnc_RTD1406 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010101111110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1406)
);
fnc_RTD1407 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010101111111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1407)
);
fnc_RTD1408 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010110000000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1408)
);
fnc_RTD1409 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010110000001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1409)
);
fnc_RTD1410 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010110000010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1410)
);
fnc_RTD1411 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010110000011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1411)
);
fnc_RTD1412 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010110000100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1412)
);
fnc_RTD1413 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010110000101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1413)
);
fnc_RTD1414 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010110000110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1414)
);
fnc_RTD1415 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010110000111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1415)
);
fnc_RTD1416 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010110001000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1416)
);
fnc_RTD1417 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010110001001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1417)
);
fnc_RTD1418 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010110001010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1418)
);
fnc_RTD1419 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010110001011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1419)
);
fnc_RTD1420 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010110001100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1420)
);
fnc_RTD1421 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010110001101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1421)
);
fnc_RTD1422 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010110001110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1422)
);
fnc_RTD1423 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010110001111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1423)
);
fnc_RTD1424 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010110010000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1424)
);
fnc_RTD1425 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010110010001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1425)
);
fnc_RTD1426 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010110010010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1426)
);
fnc_RTD1427 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010110010011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1427)
);
fnc_RTD1428 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010110010100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1428)
);
fnc_RTD1429 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010110010101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1429)
);
fnc_RTD1430 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010110010110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1430)
);
fnc_RTD1431 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010110010111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1431)
);
fnc_RTD1432 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010110011000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1432)
);
fnc_RTD1433 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010110011001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1433)
);
fnc_RTD1434 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010110011010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1434)
);
fnc_RTD1435 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010110011011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1435)
);
fnc_RTD1436 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010110011100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1436)
);
fnc_RTD1437 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010110011101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1437)
);
fnc_RTD1438 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010110011110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1438)
);
fnc_RTD1439 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010110011111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1439)
);
fnc_RTD1440 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010110100000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1440)
);
fnc_RTD1441 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010110100001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1441)
);
fnc_RTD1442 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010110100010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1442)
);
fnc_RTD1443 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010110100011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1443)
);
fnc_RTD1444 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010110100100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1444)
);
fnc_RTD1445 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010110100101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1445)
);
fnc_RTD1446 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010110100110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1446)
);
fnc_RTD1447 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010110100111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1447)
);
fnc_RTD1448 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010110101000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1448)
);
fnc_RTD1449 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010110101001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1449)
);
fnc_RTD1450 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010110101010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1450)
);
fnc_RTD1451 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010110101011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1451)
);
fnc_RTD1452 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010110101100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1452)
);
fnc_RTD1453 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010110101101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1453)
);
fnc_RTD1454 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010110101110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1454)
);
fnc_RTD1455 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010110101111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1455)
);
fnc_RTD1456 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010110110000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1456)
);
fnc_RTD1457 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010110110001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1457)
);
fnc_RTD1458 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010110110010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1458)
);
fnc_RTD1459 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010110110011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1459)
);
fnc_RTD1460 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010110110100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1460)
);
fnc_RTD1461 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010110110101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1461)
);
fnc_RTD1462 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010110110110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1462)
);
fnc_RTD1463 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010110110111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1463)
);
fnc_RTD1464 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010110111000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1464)
);
fnc_RTD1465 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010110111001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1465)
);
fnc_RTD1466 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010110111010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1466)
);
fnc_RTD1467 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010110111011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1467)
);
fnc_RTD1468 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010110111100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1468)
);
fnc_RTD1469 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010110111101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1469)
);
fnc_RTD1470 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010110111110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1470)
);
fnc_RTD1471 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010110111111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1471)
);
fnc_RTD1472 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010111000000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1472)
);
fnc_RTD1473 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010111000001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1473)
);
fnc_RTD1474 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010111000010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1474)
);
fnc_RTD1475 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010111000011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1475)
);
fnc_RTD1476 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010111000100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1476)
);
fnc_RTD1477 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010111000101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1477)
);
fnc_RTD1478 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010111000110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1478)
);
fnc_RTD1479 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010111000111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1479)
);
fnc_RTD1480 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010111001000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1480)
);
fnc_RTD1481 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010111001001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1481)
);
fnc_RTD1482 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010111001010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1482)
);
fnc_RTD1483 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010111001011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1483)
);
fnc_RTD1484 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010111001100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1484)
);
fnc_RTD1485 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010111001101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1485)
);
fnc_RTD1486 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010111001110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1486)
);
fnc_RTD1487 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010111001111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1487)
);
fnc_RTD1488 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010111010000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1488)
);
fnc_RTD1489 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010111010001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1489)
);
fnc_RTD1490 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010111010010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1490)
);
fnc_RTD1491 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010111010011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1491)
);
fnc_RTD1492 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010111010100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1492)
);
fnc_RTD1493 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010111010101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1493)
);
fnc_RTD1494 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010111010110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1494)
);
fnc_RTD1495 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010111010111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1495)
);
fnc_RTD1496 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010111011000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1496)
);
fnc_RTD1497 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010111011001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1497)
);
fnc_RTD1498 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010111011010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1498)
);
fnc_RTD1499 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010111011011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1499)
);
fnc_RTD1500 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010111011100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1500)
);
fnc_RTD1501 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010111011101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1501)
);
fnc_RTD1502 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010111011110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1502)
);
fnc_RTD1503 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010111011111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1503)
);
fnc_RTD1504 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010111100000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1504)
);
fnc_RTD1505 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010111100001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1505)
);
fnc_RTD1506 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010111100010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1506)
);
fnc_RTD1507 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010111100011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1507)
);
fnc_RTD1508 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010111100100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1508)
);
fnc_RTD1509 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010111100101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1509)
);
fnc_RTD1510 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010111100110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1510)
);
fnc_RTD1511 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010111100111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1511)
);
fnc_RTD1512 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010111101000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1512)
);
fnc_RTD1513 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010111101001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1513)
);
fnc_RTD1514 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010111101010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1514)
);
fnc_RTD1515 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010111101011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1515)
);
fnc_RTD1516 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010111101100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1516)
);
fnc_RTD1517 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010111101101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1517)
);
fnc_RTD1518 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010111101110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1518)
);
fnc_RTD1519 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010111101111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1519)
);
fnc_RTD1520 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010111110000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1520)
);
fnc_RTD1521 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010111110001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1521)
);
fnc_RTD1522 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010111110010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1522)
);
fnc_RTD1523 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010111110011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1523)
);
fnc_RTD1524 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010111110100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1524)
);
fnc_RTD1525 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010111110101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1525)
);
fnc_RTD1526 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010111110110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1526)
);
fnc_RTD1527 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010111110111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1527)
);
fnc_RTD1528 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010111111000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1528)
);
fnc_RTD1529 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010111111001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1529)
);
fnc_RTD1530 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010111111010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1530)
);
fnc_RTD1531 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010111111011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1531)
);
fnc_RTD1532 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010111111100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1532)
);
fnc_RTD1533 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010111111101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1533)
);
fnc_RTD1534 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010111111110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1534)
);
fnc_RTD1535 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010111111111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1535)
);
fnc_RTD1536 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011000000000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1536)
);
fnc_RTD1537 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011000000001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1537)
);
fnc_RTD1538 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011000000010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1538)
);
fnc_RTD1539 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011000000011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1539)
);
fnc_RTD1540 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011000000100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1540)
);
fnc_RTD1541 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011000000101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1541)
);
fnc_RTD1542 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011000000110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1542)
);
fnc_RTD1543 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011000000111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1543)
);
fnc_RTD1544 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011000001000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1544)
);
fnc_RTD1545 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011000001001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1545)
);
fnc_RTD1546 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011000001010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1546)
);
fnc_RTD1547 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011000001011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1547)
);
fnc_RTD1548 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011000001100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1548)
);
fnc_RTD1549 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011000001101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1549)
);
fnc_RTD1550 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011000001110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1550)
);
fnc_RTD1551 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011000001111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1551)
);
fnc_RTD1552 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011000010000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1552)
);
fnc_RTD1553 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011000010001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1553)
);
fnc_RTD1554 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011000010010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1554)
);
fnc_RTD1555 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011000010011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1555)
);
fnc_RTD1556 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011000010100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1556)
);
fnc_RTD1557 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011000010101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1557)
);
fnc_RTD1558 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011000010110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1558)
);
fnc_RTD1559 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011000010111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1559)
);
fnc_RTD1560 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011000011000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1560)
);
fnc_RTD1561 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011000011001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1561)
);
fnc_RTD1562 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011000011010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1562)
);
fnc_RTD1563 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011000011011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1563)
);
fnc_RTD1564 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011000011100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1564)
);
fnc_RTD1565 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011000011101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1565)
);
fnc_RTD1566 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011000011110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1566)
);
fnc_RTD1567 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011000011111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1567)
);
fnc_RTD1568 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011000100000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1568)
);
fnc_RTD1569 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011000100001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1569)
);
fnc_RTD1570 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011000100010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1570)
);
fnc_RTD1571 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011000100011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1571)
);
fnc_RTD1572 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011000100100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1572)
);
fnc_RTD1573 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011000100101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1573)
);
fnc_RTD1574 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011000100110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1574)
);
fnc_RTD1575 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011000100111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1575)
);
fnc_RTD1576 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011000101000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1576)
);
fnc_RTD1577 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011000101001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1577)
);
fnc_RTD1578 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011000101010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1578)
);
fnc_RTD1579 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011000101011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1579)
);
fnc_RTD1580 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011000101100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1580)
);
fnc_RTD1581 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011000101101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1581)
);
fnc_RTD1582 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011000101110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1582)
);
fnc_RTD1583 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011000101111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1583)
);
fnc_RTD1584 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011000110000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1584)
);
fnc_RTD1585 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011000110001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1585)
);
fnc_RTD1586 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011000110010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1586)
);
fnc_RTD1587 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011000110011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1587)
);
fnc_RTD1588 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011000110100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1588)
);
fnc_RTD1589 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011000110101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1589)
);
fnc_RTD1590 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011000110110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1590)
);
fnc_RTD1591 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011000110111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1591)
);
fnc_RTD1592 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011000111000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1592)
);
fnc_RTD1593 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011000111001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1593)
);
fnc_RTD1594 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011000111010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1594)
);
fnc_RTD1595 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011000111011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1595)
);
fnc_RTD1596 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011000111100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1596)
);
fnc_RTD1597 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011000111101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1597)
);
fnc_RTD1598 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011000111110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1598)
);
fnc_RTD1599 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011000111111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1599)
);
fnc_RTD1600 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011001000000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1600)
);
fnc_RTD1601 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011001000001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1601)
);
fnc_RTD1602 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011001000010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1602)
);
fnc_RTD1603 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011001000011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1603)
);
fnc_RTD1604 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011001000100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1604)
);
fnc_RTD1605 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011001000101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1605)
);
fnc_RTD1606 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011001000110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1606)
);
fnc_RTD1607 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011001000111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1607)
);
fnc_RTD1608 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011001001000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1608)
);
fnc_RTD1609 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011001001001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1609)
);
fnc_RTD1610 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011001001010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1610)
);
fnc_RTD1611 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011001001011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1611)
);
fnc_RTD1612 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011001001100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1612)
);
fnc_RTD1613 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011001001101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1613)
);
fnc_RTD1614 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011001001110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1614)
);
fnc_RTD1615 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011001001111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1615)
);
fnc_RTD1616 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011001010000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1616)
);
fnc_RTD1617 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011001010001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1617)
);
fnc_RTD1618 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011001010010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1618)
);
fnc_RTD1619 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011001010011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1619)
);
fnc_RTD1620 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011001010100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1620)
);
fnc_RTD1621 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011001010101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1621)
);
fnc_RTD1622 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011001010110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1622)
);
fnc_RTD1623 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011001010111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1623)
);
fnc_RTD1624 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011001011000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1624)
);
fnc_RTD1625 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011001011001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1625)
);
fnc_RTD1626 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011001011010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1626)
);
fnc_RTD1627 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011001011011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1627)
);
fnc_RTD1628 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011001011100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1628)
);
fnc_RTD1629 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011001011101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1629)
);
fnc_RTD1630 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011001011110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1630)
);
fnc_RTD1631 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011001011111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1631)
);
fnc_RTD1632 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011001100000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1632)
);
fnc_RTD1633 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011001100001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1633)
);
fnc_RTD1634 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011001100010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1634)
);
fnc_RTD1635 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011001100011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1635)
);
fnc_RTD1636 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011001100100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1636)
);
fnc_RTD1637 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011001100101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1637)
);
fnc_RTD1638 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011001100110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1638)
);
fnc_RTD1639 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011001100111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1639)
);
fnc_RTD1640 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011001101000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1640)
);
fnc_RTD1641 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011001101001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1641)
);
fnc_RTD1642 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011001101010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1642)
);
fnc_RTD1643 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011001101011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1643)
);
fnc_RTD1644 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011001101100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1644)
);
fnc_RTD1645 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011001101101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1645)
);
fnc_RTD1646 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011001101110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1646)
);
fnc_RTD1647 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011001101111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1647)
);
fnc_RTD1648 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011001110000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1648)
);
fnc_RTD1649 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011001110001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1649)
);
fnc_RTD1650 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011001110010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1650)
);
fnc_RTD1651 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011001110011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1651)
);
fnc_RTD1652 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011001110100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1652)
);
fnc_RTD1653 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011001110101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1653)
);
fnc_RTD1654 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011001110110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1654)
);
fnc_RTD1655 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011001110111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1655)
);
fnc_RTD1656 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011001111000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1656)
);
fnc_RTD1657 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011001111001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1657)
);
fnc_RTD1658 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011001111010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1658)
);
fnc_RTD1659 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011001111011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1659)
);
fnc_RTD1660 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011001111100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1660)
);
fnc_RTD1661 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011001111101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1661)
);
fnc_RTD1662 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011001111110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1662)
);
fnc_RTD1663 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011001111111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1663)
);
fnc_RTD1664 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011010000000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1664)
);
fnc_RTD1665 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011010000001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1665)
);
fnc_RTD1666 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011010000010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1666)
);
fnc_RTD1667 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011010000011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1667)
);
fnc_RTD1668 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011010000100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1668)
);
fnc_RTD1669 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011010000101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1669)
);
fnc_RTD1670 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011010000110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1670)
);
fnc_RTD1671 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011010000111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1671)
);
fnc_RTD1672 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011010001000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1672)
);
fnc_RTD1673 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011010001001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1673)
);
fnc_RTD1674 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011010001010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1674)
);
fnc_RTD1675 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011010001011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1675)
);
fnc_RTD1676 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011010001100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1676)
);
fnc_RTD1677 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011010001101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1677)
);
fnc_RTD1678 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011010001110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1678)
);
fnc_RTD1679 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011010001111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1679)
);
fnc_RTD1680 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011010010000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1680)
);
fnc_RTD1681 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011010010001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1681)
);
fnc_RTD1682 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011010010010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1682)
);
fnc_RTD1683 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011010010011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1683)
);
fnc_RTD1684 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011010010100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1684)
);
fnc_RTD1685 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011010010101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1685)
);
fnc_RTD1686 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011010010110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1686)
);
fnc_RTD1687 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011010010111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1687)
);
fnc_RTD1688 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011010011000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1688)
);
fnc_RTD1689 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011010011001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1689)
);
fnc_RTD1690 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011010011010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1690)
);
fnc_RTD1691 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011010011011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1691)
);
fnc_RTD1692 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011010011100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1692)
);
fnc_RTD1693 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011010011101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1693)
);
fnc_RTD1694 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011010011110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1694)
);
fnc_RTD1695 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011010011111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1695)
);
fnc_RTD1696 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011010100000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1696)
);
fnc_RTD1697 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011010100001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1697)
);
fnc_RTD1698 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011010100010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1698)
);
fnc_RTD1699 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011010100011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1699)
);
fnc_RTD1700 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011010100100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1700)
);
fnc_RTD1701 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011010100101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1701)
);
fnc_RTD1702 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011010100110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1702)
);
fnc_RTD1703 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011010100111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1703)
);
fnc_RTD1704 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011010101000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1704)
);
fnc_RTD1705 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011010101001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1705)
);
fnc_RTD1706 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011010101010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1706)
);
fnc_RTD1707 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011010101011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1707)
);
fnc_RTD1708 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011010101100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1708)
);
fnc_RTD1709 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011010101101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1709)
);
fnc_RTD1710 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011010101110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1710)
);
fnc_RTD1711 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011010101111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1711)
);
fnc_RTD1712 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011010110000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1712)
);
fnc_RTD1713 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011010110001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1713)
);
fnc_RTD1714 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011010110010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1714)
);
fnc_RTD1715 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011010110011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1715)
);
fnc_RTD1716 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011010110100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1716)
);
fnc_RTD1717 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011010110101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1717)
);
fnc_RTD1718 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011010110110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1718)
);
fnc_RTD1719 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011010110111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1719)
);
fnc_RTD1720 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011010111000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1720)
);
fnc_RTD1721 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011010111001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1721)
);
fnc_RTD1722 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011010111010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1722)
);
fnc_RTD1723 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011010111011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1723)
);
fnc_RTD1724 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011010111100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1724)
);
fnc_RTD1725 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011010111101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1725)
);
fnc_RTD1726 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011010111110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1726)
);
fnc_RTD1727 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011010111111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1727)
);
fnc_RTD1728 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011011000000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1728)
);
fnc_RTD1729 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011011000001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1729)
);
fnc_RTD1730 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011011000010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1730)
);
fnc_RTD1731 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011011000011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1731)
);
fnc_RTD1732 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011011000100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1732)
);
fnc_RTD1733 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011011000101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1733)
);
fnc_RTD1734 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011011000110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1734)
);
fnc_RTD1735 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011011000111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1735)
);
fnc_RTD1736 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011011001000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1736)
);
fnc_RTD1737 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011011001001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1737)
);
fnc_RTD1738 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011011001010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1738)
);
fnc_RTD1739 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011011001011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1739)
);
fnc_RTD1740 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011011001100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1740)
);
fnc_RTD1741 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011011001101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1741)
);
fnc_RTD1742 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011011001110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1742)
);
fnc_RTD1743 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011011001111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1743)
);
fnc_RTD1744 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011011010000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1744)
);
fnc_RTD1745 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011011010001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1745)
);
fnc_RTD1746 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011011010010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1746)
);
fnc_RTD1747 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011011010011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1747)
);
fnc_RTD1748 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011011010100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1748)
);
fnc_RTD1749 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011011010101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1749)
);
fnc_RTD1750 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011011010110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1750)
);
fnc_RTD1751 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011011010111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1751)
);
fnc_RTD1752 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011011011000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1752)
);
fnc_RTD1753 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011011011001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1753)
);
fnc_RTD1754 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011011011010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1754)
);
fnc_RTD1755 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011011011011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1755)
);
fnc_RTD1756 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011011011100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1756)
);
fnc_RTD1757 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011011011101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1757)
);
fnc_RTD1758 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011011011110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1758)
);
fnc_RTD1759 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011011011111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1759)
);
fnc_RTD1760 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011011100000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1760)
);
fnc_RTD1761 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011011100001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1761)
);
fnc_RTD1762 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011011100010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1762)
);
fnc_RTD1763 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011011100011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1763)
);
fnc_RTD1764 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011011100100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1764)
);
fnc_RTD1765 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011011100101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1765)
);
fnc_RTD1766 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011011100110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1766)
);
fnc_RTD1767 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011011100111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1767)
);
fnc_RTD1768 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011011101000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1768)
);
fnc_RTD1769 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011011101001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1769)
);
fnc_RTD1770 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011011101010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1770)
);
fnc_RTD1771 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011011101011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1771)
);
fnc_RTD1772 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011011101100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1772)
);
fnc_RTD1773 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011011101101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1773)
);
fnc_RTD1774 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011011101110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1774)
);
fnc_RTD1775 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011011101111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1775)
);
fnc_RTD1776 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011011110000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1776)
);
fnc_RTD1777 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011011110001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1777)
);
fnc_RTD1778 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011011110010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1778)
);
fnc_RTD1779 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011011110011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1779)
);
fnc_RTD1780 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011011110100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1780)
);
fnc_RTD1781 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011011110101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1781)
);
fnc_RTD1782 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011011110110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1782)
);
fnc_RTD1783 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011011110111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1783)
);
fnc_RTD1784 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011011111000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1784)
);
fnc_RTD1785 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011011111001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1785)
);
fnc_RTD1786 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011011111010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1786)
);
fnc_RTD1787 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011011111011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1787)
);
fnc_RTD1788 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011011111100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1788)
);
fnc_RTD1789 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011011111101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1789)
);
fnc_RTD1790 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011011111110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1790)
);
fnc_RTD1791 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011011111111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1791)
);
fnc_RTD1792 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011100000000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1792)
);
fnc_RTD1793 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011100000001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1793)
);
fnc_RTD1794 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011100000010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1794)
);
fnc_RTD1795 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011100000011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1795)
);
fnc_RTD1796 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011100000100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1796)
);
fnc_RTD1797 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011100000101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1797)
);
fnc_RTD1798 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011100000110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1798)
);
fnc_RTD1799 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011100000111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1799)
);
fnc_RTD1800 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011100001000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1800)
);
fnc_RTD1801 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011100001001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1801)
);
fnc_RTD1802 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011100001010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1802)
);
fnc_RTD1803 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011100001011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1803)
);
fnc_RTD1804 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011100001100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1804)
);
fnc_RTD1805 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011100001101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1805)
);
fnc_RTD1806 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011100001110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1806)
);
fnc_RTD1807 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011100001111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1807)
);
fnc_RTD1808 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011100010000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1808)
);
fnc_RTD1809 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011100010001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1809)
);
fnc_RTD1810 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011100010010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1810)
);
fnc_RTD1811 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011100010011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1811)
);
fnc_RTD1812 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011100010100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1812)
);
fnc_RTD1813 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011100010101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1813)
);
fnc_RTD1814 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011100010110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1814)
);
fnc_RTD1815 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011100010111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1815)
);
fnc_RTD1816 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011100011000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1816)
);
fnc_RTD1817 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011100011001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1817)
);
fnc_RTD1818 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011100011010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1818)
);
fnc_RTD1819 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011100011011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1819)
);
fnc_RTD1820 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011100011100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1820)
);
fnc_RTD1821 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011100011101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1821)
);
fnc_RTD1822 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011100011110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1822)
);
fnc_RTD1823 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011100011111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1823)
);
fnc_RTD1824 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011100100000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1824)
);
fnc_RTD1825 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011100100001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1825)
);
fnc_RTD1826 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011100100010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1826)
);
fnc_RTD1827 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011100100011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1827)
);
fnc_RTD1828 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011100100100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1828)
);
fnc_RTD1829 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011100100101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1829)
);
fnc_RTD1830 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011100100110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1830)
);
fnc_RTD1831 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011100100111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1831)
);
fnc_RTD1832 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011100101000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1832)
);
fnc_RTD1833 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011100101001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1833)
);
fnc_RTD1834 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011100101010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1834)
);
fnc_RTD1835 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011100101011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1835)
);
fnc_RTD1836 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011100101100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1836)
);
fnc_RTD1837 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011100101101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1837)
);
fnc_RTD1838 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011100101110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1838)
);
fnc_RTD1839 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011100101111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1839)
);
fnc_RTD1840 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011100110000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1840)
);
fnc_RTD1841 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011100110001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1841)
);
fnc_RTD1842 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011100110010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1842)
);
fnc_RTD1843 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011100110011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1843)
);
fnc_RTD1844 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011100110100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1844)
);
fnc_RTD1845 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011100110101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1845)
);
fnc_RTD1846 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011100110110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1846)
);
fnc_RTD1847 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011100110111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1847)
);
fnc_RTD1848 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011100111000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1848)
);
fnc_RTD1849 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011100111001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1849)
);
fnc_RTD1850 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011100111010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1850)
);
fnc_RTD1851 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011100111011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1851)
);
fnc_RTD1852 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011100111100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1852)
);
fnc_RTD1853 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011100111101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1853)
);
fnc_RTD1854 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011100111110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1854)
);
fnc_RTD1855 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011100111111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1855)
);
fnc_RTD1856 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011101000000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1856)
);
fnc_RTD1857 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011101000001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1857)
);
fnc_RTD1858 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011101000010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1858)
);
fnc_RTD1859 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011101000011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1859)
);
fnc_RTD1860 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011101000100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1860)
);
fnc_RTD1861 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011101000101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1861)
);
fnc_RTD1862 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011101000110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1862)
);
fnc_RTD1863 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011101000111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1863)
);
fnc_RTD1864 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011101001000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1864)
);
fnc_RTD1865 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011101001001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1865)
);
fnc_RTD1866 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011101001010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1866)
);
fnc_RTD1867 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011101001011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1867)
);
fnc_RTD1868 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011101001100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1868)
);
fnc_RTD1869 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011101001101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1869)
);
fnc_RTD1870 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011101001110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1870)
);
fnc_RTD1871 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011101001111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1871)
);
fnc_RTD1872 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011101010000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1872)
);
fnc_RTD1873 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011101010001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1873)
);
fnc_RTD1874 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011101010010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1874)
);
fnc_RTD1875 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011101010011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1875)
);
fnc_RTD1876 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011101010100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1876)
);
fnc_RTD1877 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011101010101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1877)
);
fnc_RTD1878 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011101010110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1878)
);
fnc_RTD1879 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011101010111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1879)
);
fnc_RTD1880 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011101011000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1880)
);
fnc_RTD1881 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011101011001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1881)
);
fnc_RTD1882 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011101011010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1882)
);
fnc_RTD1883 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011101011011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1883)
);
fnc_RTD1884 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011101011100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1884)
);
fnc_RTD1885 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011101011101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1885)
);
fnc_RTD1886 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011101011110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1886)
);
fnc_RTD1887 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011101011111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1887)
);
fnc_RTD1888 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011101100000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1888)
);
fnc_RTD1889 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011101100001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1889)
);
fnc_RTD1890 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011101100010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1890)
);
fnc_RTD1891 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011101100011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1891)
);
fnc_RTD1892 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011101100100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1892)
);
fnc_RTD1893 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011101100101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1893)
);
fnc_RTD1894 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011101100110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1894)
);
fnc_RTD1895 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011101100111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1895)
);
fnc_RTD1896 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011101101000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1896)
);
fnc_RTD1897 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011101101001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1897)
);
fnc_RTD1898 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011101101010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1898)
);
fnc_RTD1899 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011101101011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1899)
);
fnc_RTD1900 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011101101100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1900)
);
fnc_RTD1901 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011101101101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1901)
);
fnc_RTD1902 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011101101110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1902)
);
fnc_RTD1903 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011101101111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1903)
);
fnc_RTD1904 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011101110000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1904)
);
fnc_RTD1905 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011101110001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1905)
);
fnc_RTD1906 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011101110010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1906)
);
fnc_RTD1907 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011101110011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1907)
);
fnc_RTD1908 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011101110100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1908)
);
fnc_RTD1909 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011101110101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1909)
);
fnc_RTD1910 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011101110110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1910)
);
fnc_RTD1911 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011101110111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1911)
);
fnc_RTD1912 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011101111000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1912)
);
fnc_RTD1913 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011101111001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1913)
);
fnc_RTD1914 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011101111010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1914)
);
fnc_RTD1915 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011101111011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1915)
);
fnc_RTD1916 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011101111100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1916)
);
fnc_RTD1917 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011101111101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1917)
);
fnc_RTD1918 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011101111110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1918)
);
fnc_RTD1919 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011101111111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1919)
);
fnc_RTD1920 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011110000000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1920)
);
fnc_RTD1921 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011110000001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1921)
);
fnc_RTD1922 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011110000010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1922)
);
fnc_RTD1923 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011110000011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1923)
);
fnc_RTD1924 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011110000100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1924)
);
fnc_RTD1925 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011110000101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1925)
);
fnc_RTD1926 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011110000110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1926)
);
fnc_RTD1927 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011110000111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1927)
);
fnc_RTD1928 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011110001000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1928)
);
fnc_RTD1929 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011110001001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1929)
);
fnc_RTD1930 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011110001010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1930)
);
fnc_RTD1931 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011110001011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1931)
);
fnc_RTD1932 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011110001100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1932)
);
fnc_RTD1933 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011110001101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1933)
);
fnc_RTD1934 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011110001110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1934)
);
fnc_RTD1935 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011110001111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1935)
);
fnc_RTD1936 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011110010000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1936)
);
fnc_RTD1937 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011110010001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1937)
);
fnc_RTD1938 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011110010010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1938)
);
fnc_RTD1939 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011110010011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1939)
);
fnc_RTD1940 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011110010100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1940)
);
fnc_RTD1941 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011110010101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1941)
);
fnc_RTD1942 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011110010110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1942)
);
fnc_RTD1943 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011110010111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1943)
);
fnc_RTD1944 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011110011000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1944)
);
fnc_RTD1945 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011110011001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1945)
);
fnc_RTD1946 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011110011010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1946)
);
fnc_RTD1947 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011110011011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1947)
);
fnc_RTD1948 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011110011100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1948)
);
fnc_RTD1949 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011110011101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1949)
);
fnc_RTD1950 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011110011110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1950)
);
fnc_RTD1951 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011110011111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1951)
);
fnc_RTD1952 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011110100000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1952)
);
fnc_RTD1953 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011110100001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1953)
);
fnc_RTD1954 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011110100010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1954)
);
fnc_RTD1955 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011110100011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1955)
);
fnc_RTD1956 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011110100100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1956)
);
fnc_RTD1957 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011110100101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1957)
);
fnc_RTD1958 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011110100110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1958)
);
fnc_RTD1959 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011110100111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1959)
);
fnc_RTD1960 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011110101000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1960)
);
fnc_RTD1961 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011110101001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1961)
);
fnc_RTD1962 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011110101010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1962)
);
fnc_RTD1963 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011110101011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1963)
);
fnc_RTD1964 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011110101100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1964)
);
fnc_RTD1965 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011110101101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1965)
);
fnc_RTD1966 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011110101110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1966)
);
fnc_RTD1967 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011110101111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1967)
);
fnc_RTD1968 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011110110000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1968)
);
fnc_RTD1969 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011110110001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1969)
);
fnc_RTD1970 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011110110010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1970)
);
fnc_RTD1971 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011110110011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1971)
);
fnc_RTD1972 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011110110100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1972)
);
fnc_RTD1973 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011110110101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1973)
);
fnc_RTD1974 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011110110110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1974)
);
fnc_RTD1975 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011110110111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1975)
);
fnc_RTD1976 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011110111000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1976)
);
fnc_RTD1977 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011110111001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1977)
);
fnc_RTD1978 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011110111010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1978)
);
fnc_RTD1979 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011110111011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1979)
);
fnc_RTD1980 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011110111100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1980)
);
fnc_RTD1981 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011110111101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1981)
);
fnc_RTD1982 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011110111110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1982)
);
fnc_RTD1983 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011110111111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1983)
);
fnc_RTD1984 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011111000000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1984)
);
fnc_RTD1985 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011111000001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1985)
);
fnc_RTD1986 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011111000010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1986)
);
fnc_RTD1987 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011111000011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1987)
);
fnc_RTD1988 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011111000100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1988)
);
fnc_RTD1989 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011111000101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1989)
);
fnc_RTD1990 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011111000110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1990)
);
fnc_RTD1991 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011111000111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1991)
);
fnc_RTD1992 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011111001000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1992)
);
fnc_RTD1993 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011111001001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1993)
);
fnc_RTD1994 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011111001010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1994)
);
fnc_RTD1995 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011111001011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1995)
);
fnc_RTD1996 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011111001100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1996)
);
fnc_RTD1997 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011111001101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1997)
);
fnc_RTD1998 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011111001110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1998)
);
fnc_RTD1999 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011111001111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(1999)
);
fnc_RTD2000 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011111010000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2000)
);
fnc_RTD2001 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011111010001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2001)
);
fnc_RTD2002 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011111010010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2002)
);
fnc_RTD2003 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011111010011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2003)
);
fnc_RTD2004 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011111010100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2004)
);
fnc_RTD2005 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011111010101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2005)
);
fnc_RTD2006 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011111010110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2006)
);
fnc_RTD2007 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011111010111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2007)
);
fnc_RTD2008 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011111011000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2008)
);
fnc_RTD2009 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011111011001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2009)
);
fnc_RTD2010 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011111011010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2010)
);
fnc_RTD2011 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011111011011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2011)
);
fnc_RTD2012 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011111011100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2012)
);
fnc_RTD2013 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011111011101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2013)
);
fnc_RTD2014 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011111011110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2014)
);
fnc_RTD2015 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011111011111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2015)
);
fnc_RTD2016 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011111100000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2016)
);
fnc_RTD2017 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011111100001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2017)
);
fnc_RTD2018 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011111100010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2018)
);
fnc_RTD2019 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011111100011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2019)
);
fnc_RTD2020 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011111100100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2020)
);
fnc_RTD2021 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011111100101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2021)
);
fnc_RTD2022 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011111100110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2022)
);
fnc_RTD2023 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011111100111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2023)
);
fnc_RTD2024 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011111101000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2024)
);
fnc_RTD2025 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011111101001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2025)
);
fnc_RTD2026 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011111101010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2026)
);
fnc_RTD2027 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011111101011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2027)
);
fnc_RTD2028 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011111101100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2028)
);
fnc_RTD2029 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011111101101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2029)
);
fnc_RTD2030 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011111101110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2030)
);
fnc_RTD2031 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011111101111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2031)
);
fnc_RTD2032 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011111110000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2032)
);
fnc_RTD2033 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011111110001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2033)
);
fnc_RTD2034 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011111110010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2034)
);
fnc_RTD2035 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011111110011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2035)
);
fnc_RTD2036 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011111110100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2036)
);
fnc_RTD2037 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011111110101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2037)
);
fnc_RTD2038 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011111110110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2038)
);
fnc_RTD2039 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011111110111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2039)
);
fnc_RTD2040 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011111111000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2040)
);
fnc_RTD2041 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011111111001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2041)
);
fnc_RTD2042 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011111111010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2042)
);
fnc_RTD2043 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011111111011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2043)
);
fnc_RTD2044 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011111111100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2044)
);
fnc_RTD2045 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011111111101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2045)
);
fnc_RTD2046 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011111111110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2046)
);
fnc_RTD2047 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000011111111111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2047)
);
fnc_RTD2048 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100000000000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2048)
);
fnc_RTD2049 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100000000001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2049)
);
fnc_RTD2050 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100000000010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2050)
);
fnc_RTD2051 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100000000011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2051)
);
fnc_RTD2052 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100000000100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2052)
);
fnc_RTD2053 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100000000101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2053)
);
fnc_RTD2054 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100000000110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2054)
);
fnc_RTD2055 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100000000111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2055)
);
fnc_RTD2056 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100000001000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2056)
);
fnc_RTD2057 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100000001001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2057)
);
fnc_RTD2058 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100000001010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2058)
);
fnc_RTD2059 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100000001011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2059)
);
fnc_RTD2060 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100000001100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2060)
);
fnc_RTD2061 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100000001101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2061)
);
fnc_RTD2062 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100000001110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2062)
);
fnc_RTD2063 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100000001111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2063)
);
fnc_RTD2064 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100000010000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2064)
);
fnc_RTD2065 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100000010001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2065)
);
fnc_RTD2066 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100000010010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2066)
);
fnc_RTD2067 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100000010011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2067)
);
fnc_RTD2068 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100000010100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2068)
);
fnc_RTD2069 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100000010101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2069)
);
fnc_RTD2070 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100000010110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2070)
);
fnc_RTD2071 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100000010111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2071)
);
fnc_RTD2072 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100000011000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2072)
);
fnc_RTD2073 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100000011001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2073)
);
fnc_RTD2074 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100000011010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2074)
);
fnc_RTD2075 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100000011011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2075)
);
fnc_RTD2076 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100000011100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2076)
);
fnc_RTD2077 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100000011101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2077)
);
fnc_RTD2078 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100000011110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2078)
);
fnc_RTD2079 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100000011111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2079)
);
fnc_RTD2080 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100000100000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2080)
);
fnc_RTD2081 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100000100001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2081)
);
fnc_RTD2082 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100000100010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2082)
);
fnc_RTD2083 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100000100011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2083)
);
fnc_RTD2084 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100000100100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2084)
);
fnc_RTD2085 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100000100101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2085)
);
fnc_RTD2086 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100000100110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2086)
);
fnc_RTD2087 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100000100111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2087)
);
fnc_RTD2088 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100000101000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2088)
);
fnc_RTD2089 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100000101001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2089)
);
fnc_RTD2090 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100000101010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2090)
);
fnc_RTD2091 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100000101011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2091)
);
fnc_RTD2092 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100000101100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2092)
);
fnc_RTD2093 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100000101101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2093)
);
fnc_RTD2094 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100000101110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2094)
);
fnc_RTD2095 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100000101111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2095)
);
fnc_RTD2096 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100000110000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2096)
);
fnc_RTD2097 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100000110001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2097)
);
fnc_RTD2098 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100000110010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2098)
);
fnc_RTD2099 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100000110011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2099)
);
fnc_RTD2100 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100000110100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2100)
);
fnc_RTD2101 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100000110101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2101)
);
fnc_RTD2102 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100000110110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2102)
);
fnc_RTD2103 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100000110111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2103)
);
fnc_RTD2104 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100000111000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2104)
);
fnc_RTD2105 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100000111001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2105)
);
fnc_RTD2106 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100000111010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2106)
);
fnc_RTD2107 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100000111011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2107)
);
fnc_RTD2108 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100000111100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2108)
);
fnc_RTD2109 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100000111101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2109)
);
fnc_RTD2110 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100000111110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2110)
);
fnc_RTD2111 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100000111111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2111)
);
fnc_RTD2112 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100001000000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2112)
);
fnc_RTD2113 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100001000001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2113)
);
fnc_RTD2114 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100001000010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2114)
);
fnc_RTD2115 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100001000011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2115)
);
fnc_RTD2116 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100001000100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2116)
);
fnc_RTD2117 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100001000101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2117)
);
fnc_RTD2118 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100001000110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2118)
);
fnc_RTD2119 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100001000111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2119)
);
fnc_RTD2120 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100001001000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2120)
);
fnc_RTD2121 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100001001001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2121)
);
fnc_RTD2122 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100001001010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2122)
);
fnc_RTD2123 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100001001011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2123)
);
fnc_RTD2124 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100001001100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2124)
);
fnc_RTD2125 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100001001101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2125)
);
fnc_RTD2126 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100001001110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2126)
);
fnc_RTD2127 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100001001111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2127)
);
fnc_RTD2128 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100001010000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2128)
);
fnc_RTD2129 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100001010001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2129)
);
fnc_RTD2130 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100001010010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2130)
);
fnc_RTD2131 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100001010011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2131)
);
fnc_RTD2132 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100001010100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2132)
);
fnc_RTD2133 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100001010101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2133)
);
fnc_RTD2134 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100001010110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2134)
);
fnc_RTD2135 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100001010111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2135)
);
fnc_RTD2136 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100001011000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2136)
);
fnc_RTD2137 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100001011001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2137)
);
fnc_RTD2138 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100001011010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2138)
);
fnc_RTD2139 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100001011011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2139)
);
fnc_RTD2140 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100001011100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2140)
);
fnc_RTD2141 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100001011101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2141)
);
fnc_RTD2142 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100001011110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2142)
);
fnc_RTD2143 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100001011111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2143)
);
fnc_RTD2144 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100001100000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2144)
);
fnc_RTD2145 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100001100001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2145)
);
fnc_RTD2146 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100001100010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2146)
);
fnc_RTD2147 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100001100011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2147)
);
fnc_RTD2148 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100001100100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2148)
);
fnc_RTD2149 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100001100101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2149)
);
fnc_RTD2150 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100001100110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2150)
);
fnc_RTD2151 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100001100111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2151)
);
fnc_RTD2152 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100001101000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2152)
);
fnc_RTD2153 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100001101001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2153)
);
fnc_RTD2154 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100001101010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2154)
);
fnc_RTD2155 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100001101011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2155)
);
fnc_RTD2156 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100001101100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2156)
);
fnc_RTD2157 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100001101101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2157)
);
fnc_RTD2158 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100001101110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2158)
);
fnc_RTD2159 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100001101111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2159)
);
fnc_RTD2160 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100001110000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2160)
);
fnc_RTD2161 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100001110001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2161)
);
fnc_RTD2162 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100001110010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2162)
);
fnc_RTD2163 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100001110011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2163)
);
fnc_RTD2164 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100001110100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2164)
);
fnc_RTD2165 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100001110101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2165)
);
fnc_RTD2166 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100001110110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2166)
);
fnc_RTD2167 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100001110111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2167)
);
fnc_RTD2168 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100001111000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2168)
);
fnc_RTD2169 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100001111001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2169)
);
fnc_RTD2170 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100001111010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2170)
);
fnc_RTD2171 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100001111011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2171)
);
fnc_RTD2172 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100001111100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2172)
);
fnc_RTD2173 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100001111101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2173)
);
fnc_RTD2174 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100001111110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2174)
);
fnc_RTD2175 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100001111111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2175)
);
fnc_RTD2176 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100010000000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2176)
);
fnc_RTD2177 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100010000001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2177)
);
fnc_RTD2178 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100010000010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2178)
);
fnc_RTD2179 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100010000011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2179)
);
fnc_RTD2180 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100010000100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2180)
);
fnc_RTD2181 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100010000101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2181)
);
fnc_RTD2182 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100010000110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2182)
);
fnc_RTD2183 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100010000111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2183)
);
fnc_RTD2184 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100010001000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2184)
);
fnc_RTD2185 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100010001001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2185)
);
fnc_RTD2186 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100010001010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2186)
);
fnc_RTD2187 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100010001011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2187)
);
fnc_RTD2188 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100010001100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2188)
);
fnc_RTD2189 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100010001101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2189)
);
fnc_RTD2190 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100010001110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2190)
);
fnc_RTD2191 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100010001111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2191)
);
fnc_RTD2192 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100010010000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2192)
);
fnc_RTD2193 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100010010001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2193)
);
fnc_RTD2194 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100010010010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2194)
);
fnc_RTD2195 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100010010011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2195)
);
fnc_RTD2196 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100010010100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2196)
);
fnc_RTD2197 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100010010101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2197)
);
fnc_RTD2198 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100010010110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2198)
);
fnc_RTD2199 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100010010111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2199)
);
fnc_RTD2200 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100010011000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2200)
);
fnc_RTD2201 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100010011001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2201)
);
fnc_RTD2202 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100010011010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2202)
);
fnc_RTD2203 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100010011011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2203)
);
fnc_RTD2204 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100010011100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2204)
);
fnc_RTD2205 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100010011101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2205)
);
fnc_RTD2206 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100010011110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2206)
);
fnc_RTD2207 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100010011111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2207)
);
fnc_RTD2208 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100010100000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2208)
);
fnc_RTD2209 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100010100001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2209)
);
fnc_RTD2210 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100010100010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2210)
);
fnc_RTD2211 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100010100011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2211)
);
fnc_RTD2212 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100010100100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2212)
);
fnc_RTD2213 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100010100101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2213)
);
fnc_RTD2214 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100010100110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2214)
);
fnc_RTD2215 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100010100111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2215)
);
fnc_RTD2216 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100010101000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2216)
);
fnc_RTD2217 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100010101001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2217)
);
fnc_RTD2218 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100010101010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2218)
);
fnc_RTD2219 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100010101011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2219)
);
fnc_RTD2220 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100010101100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2220)
);
fnc_RTD2221 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100010101101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2221)
);
fnc_RTD2222 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100010101110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2222)
);
fnc_RTD2223 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100010101111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2223)
);
fnc_RTD2224 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100010110000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2224)
);
fnc_RTD2225 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100010110001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2225)
);
fnc_RTD2226 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100010110010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2226)
);
fnc_RTD2227 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100010110011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2227)
);
fnc_RTD2228 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100010110100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2228)
);
fnc_RTD2229 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100010110101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2229)
);
fnc_RTD2230 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100010110110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2230)
);
fnc_RTD2231 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100010110111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2231)
);
fnc_RTD2232 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100010111000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2232)
);
fnc_RTD2233 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100010111001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2233)
);
fnc_RTD2234 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100010111010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2234)
);
fnc_RTD2235 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100010111011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2235)
);
fnc_RTD2236 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100010111100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2236)
);
fnc_RTD2237 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100010111101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2237)
);
fnc_RTD2238 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100010111110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2238)
);
fnc_RTD2239 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100010111111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2239)
);
fnc_RTD2240 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100011000000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2240)
);
fnc_RTD2241 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100011000001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2241)
);
fnc_RTD2242 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100011000010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2242)
);
fnc_RTD2243 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100011000011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2243)
);
fnc_RTD2244 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100011000100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2244)
);
fnc_RTD2245 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100011000101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2245)
);
fnc_RTD2246 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100011000110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2246)
);
fnc_RTD2247 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100011000111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2247)
);
fnc_RTD2248 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100011001000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2248)
);
fnc_RTD2249 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100011001001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2249)
);
fnc_RTD2250 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100011001010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2250)
);
fnc_RTD2251 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100011001011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2251)
);
fnc_RTD2252 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100011001100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2252)
);
fnc_RTD2253 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100011001101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2253)
);
fnc_RTD2254 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100011001110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2254)
);
fnc_RTD2255 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100011001111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2255)
);
fnc_RTD2256 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100011010000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2256)
);
fnc_RTD2257 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100011010001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2257)
);
fnc_RTD2258 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100011010010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2258)
);
fnc_RTD2259 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100011010011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2259)
);
fnc_RTD2260 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100011010100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2260)
);
fnc_RTD2261 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100011010101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2261)
);
fnc_RTD2262 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100011010110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2262)
);
fnc_RTD2263 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100011010111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2263)
);
fnc_RTD2264 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100011011000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2264)
);
fnc_RTD2265 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100011011001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2265)
);
fnc_RTD2266 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100011011010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2266)
);
fnc_RTD2267 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100011011011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2267)
);
fnc_RTD2268 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100011011100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2268)
);
fnc_RTD2269 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100011011101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2269)
);
fnc_RTD2270 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100011011110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2270)
);
fnc_RTD2271 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100011011111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2271)
);
fnc_RTD2272 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100011100000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2272)
);
fnc_RTD2273 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100011100001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2273)
);
fnc_RTD2274 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100011100010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2274)
);
fnc_RTD2275 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100011100011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2275)
);
fnc_RTD2276 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100011100100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2276)
);
fnc_RTD2277 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100011100101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2277)
);
fnc_RTD2278 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100011100110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2278)
);
fnc_RTD2279 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100011100111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2279)
);
fnc_RTD2280 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100011101000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2280)
);
fnc_RTD2281 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100011101001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2281)
);
fnc_RTD2282 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100011101010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2282)
);
fnc_RTD2283 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100011101011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2283)
);
fnc_RTD2284 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100011101100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2284)
);
fnc_RTD2285 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100011101101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2285)
);
fnc_RTD2286 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100011101110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2286)
);
fnc_RTD2287 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100011101111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2287)
);
fnc_RTD2288 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100011110000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2288)
);
fnc_RTD2289 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100011110001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2289)
);
fnc_RTD2290 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100011110010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2290)
);
fnc_RTD2291 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100011110011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2291)
);
fnc_RTD2292 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100011110100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2292)
);
fnc_RTD2293 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100011110101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2293)
);
fnc_RTD2294 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100011110110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2294)
);
fnc_RTD2295 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100011110111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2295)
);
fnc_RTD2296 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100011111000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2296)
);
fnc_RTD2297 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100011111001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2297)
);
fnc_RTD2298 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100011111010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2298)
);
fnc_RTD2299 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100011111011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2299)
);
fnc_RTD2300 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100011111100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2300)
);
fnc_RTD2301 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100011111101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2301)
);
fnc_RTD2302 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100011111110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2302)
);
fnc_RTD2303 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100011111111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2303)
);
fnc_RTD2304 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100100000000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2304)
);
fnc_RTD2305 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100100000001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2305)
);
fnc_RTD2306 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100100000010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2306)
);
fnc_RTD2307 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100100000011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2307)
);
fnc_RTD2308 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100100000100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2308)
);
fnc_RTD2309 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100100000101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2309)
);
fnc_RTD2310 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100100000110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2310)
);
fnc_RTD2311 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100100000111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2311)
);
fnc_RTD2312 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100100001000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2312)
);
fnc_RTD2313 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100100001001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2313)
);
fnc_RTD2314 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100100001010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2314)
);
fnc_RTD2315 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100100001011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2315)
);
fnc_RTD2316 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100100001100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2316)
);
fnc_RTD2317 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100100001101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2317)
);
fnc_RTD2318 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100100001110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2318)
);
fnc_RTD2319 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100100001111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2319)
);
fnc_RTD2320 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100100010000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2320)
);
fnc_RTD2321 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100100010001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2321)
);
fnc_RTD2322 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100100010010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2322)
);
fnc_RTD2323 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100100010011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2323)
);
fnc_RTD2324 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100100010100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2324)
);
fnc_RTD2325 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100100010101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2325)
);
fnc_RTD2326 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100100010110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2326)
);
fnc_RTD2327 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100100010111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2327)
);
fnc_RTD2328 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100100011000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2328)
);
fnc_RTD2329 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100100011001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2329)
);
fnc_RTD2330 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100100011010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2330)
);
fnc_RTD2331 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100100011011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2331)
);
fnc_RTD2332 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100100011100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2332)
);
fnc_RTD2333 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100100011101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2333)
);
fnc_RTD2334 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100100011110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2334)
);
fnc_RTD2335 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100100011111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2335)
);
fnc_RTD2336 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100100100000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2336)
);
fnc_RTD2337 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100100100001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2337)
);
fnc_RTD2338 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100100100010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2338)
);
fnc_RTD2339 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100100100011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2339)
);
fnc_RTD2340 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100100100100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2340)
);
fnc_RTD2341 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100100100101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2341)
);
fnc_RTD2342 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100100100110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2342)
);
fnc_RTD2343 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100100100111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2343)
);
fnc_RTD2344 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100100101000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2344)
);
fnc_RTD2345 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100100101001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2345)
);
fnc_RTD2346 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100100101010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2346)
);
fnc_RTD2347 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100100101011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2347)
);
fnc_RTD2348 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100100101100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2348)
);
fnc_RTD2349 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100100101101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2349)
);
fnc_RTD2350 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100100101110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2350)
);
fnc_RTD2351 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100100101111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2351)
);
fnc_RTD2352 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100100110000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2352)
);
fnc_RTD2353 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100100110001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2353)
);
fnc_RTD2354 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100100110010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2354)
);
fnc_RTD2355 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100100110011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2355)
);
fnc_RTD2356 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100100110100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2356)
);
fnc_RTD2357 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100100110101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2357)
);
fnc_RTD2358 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100100110110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2358)
);
fnc_RTD2359 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100100110111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2359)
);
fnc_RTD2360 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100100111000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2360)
);
fnc_RTD2361 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100100111001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2361)
);
fnc_RTD2362 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100100111010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2362)
);
fnc_RTD2363 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100100111011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2363)
);
fnc_RTD2364 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100100111100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2364)
);
fnc_RTD2365 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100100111101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2365)
);
fnc_RTD2366 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100100111110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2366)
);
fnc_RTD2367 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100100111111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2367)
);
fnc_RTD2368 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100101000000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2368)
);
fnc_RTD2369 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100101000001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2369)
);
fnc_RTD2370 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100101000010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2370)
);
fnc_RTD2371 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100101000011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2371)
);
fnc_RTD2372 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100101000100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2372)
);
fnc_RTD2373 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100101000101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2373)
);
fnc_RTD2374 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100101000110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2374)
);
fnc_RTD2375 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100101000111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2375)
);
fnc_RTD2376 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100101001000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2376)
);
fnc_RTD2377 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100101001001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2377)
);
fnc_RTD2378 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100101001010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2378)
);
fnc_RTD2379 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100101001011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2379)
);
fnc_RTD2380 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100101001100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2380)
);
fnc_RTD2381 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100101001101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2381)
);
fnc_RTD2382 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100101001110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2382)
);
fnc_RTD2383 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100101001111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2383)
);
fnc_RTD2384 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100101010000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2384)
);
fnc_RTD2385 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100101010001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2385)
);
fnc_RTD2386 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100101010010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2386)
);
fnc_RTD2387 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100101010011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2387)
);
fnc_RTD2388 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100101010100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2388)
);
fnc_RTD2389 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100101010101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2389)
);
fnc_RTD2390 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100101010110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2390)
);
fnc_RTD2391 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100101010111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2391)
);
fnc_RTD2392 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100101011000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2392)
);
fnc_RTD2393 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100101011001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2393)
);
fnc_RTD2394 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100101011010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2394)
);
fnc_RTD2395 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100101011011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2395)
);
fnc_RTD2396 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100101011100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2396)
);
fnc_RTD2397 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100101011101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2397)
);
fnc_RTD2398 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100101011110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2398)
);
fnc_RTD2399 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100101011111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2399)
);
fnc_RTD2400 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100101100000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2400)
);
fnc_RTD2401 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100101100001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2401)
);
fnc_RTD2402 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100101100010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2402)
);
fnc_RTD2403 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100101100011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2403)
);
fnc_RTD2404 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100101100100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2404)
);
fnc_RTD2405 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100101100101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2405)
);
fnc_RTD2406 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100101100110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2406)
);
fnc_RTD2407 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100101100111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2407)
);
fnc_RTD2408 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100101101000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2408)
);
fnc_RTD2409 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100101101001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2409)
);
fnc_RTD2410 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100101101010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2410)
);
fnc_RTD2411 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100101101011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2411)
);
fnc_RTD2412 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100101101100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2412)
);
fnc_RTD2413 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100101101101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2413)
);
fnc_RTD2414 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100101101110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2414)
);
fnc_RTD2415 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100101101111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2415)
);
fnc_RTD2416 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100101110000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2416)
);
fnc_RTD2417 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100101110001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2417)
);
fnc_RTD2418 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100101110010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2418)
);
fnc_RTD2419 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100101110011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2419)
);
fnc_RTD2420 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100101110100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2420)
);
fnc_RTD2421 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100101110101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2421)
);
fnc_RTD2422 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100101110110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2422)
);
fnc_RTD2423 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100101110111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2423)
);
fnc_RTD2424 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100101111000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2424)
);
fnc_RTD2425 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100101111001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2425)
);
fnc_RTD2426 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100101111010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2426)
);
fnc_RTD2427 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100101111011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2427)
);
fnc_RTD2428 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100101111100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2428)
);
fnc_RTD2429 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100101111101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2429)
);
fnc_RTD2430 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100101111110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2430)
);
fnc_RTD2431 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100101111111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2431)
);
fnc_RTD2432 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100110000000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2432)
);
fnc_RTD2433 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100110000001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2433)
);
fnc_RTD2434 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100110000010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2434)
);
fnc_RTD2435 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100110000011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2435)
);
fnc_RTD2436 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100110000100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2436)
);
fnc_RTD2437 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100110000101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2437)
);
fnc_RTD2438 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100110000110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2438)
);
fnc_RTD2439 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100110000111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2439)
);
fnc_RTD2440 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100110001000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2440)
);
fnc_RTD2441 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100110001001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2441)
);
fnc_RTD2442 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100110001010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2442)
);
fnc_RTD2443 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100110001011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2443)
);
fnc_RTD2444 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100110001100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2444)
);
fnc_RTD2445 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100110001101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2445)
);
fnc_RTD2446 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100110001110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2446)
);
fnc_RTD2447 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100110001111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2447)
);
fnc_RTD2448 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100110010000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2448)
);
fnc_RTD2449 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100110010001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2449)
);
fnc_RTD2450 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100110010010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2450)
);
fnc_RTD2451 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100110010011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2451)
);
fnc_RTD2452 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100110010100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2452)
);
fnc_RTD2453 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100110010101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2453)
);
fnc_RTD2454 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100110010110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2454)
);
fnc_RTD2455 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100110010111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2455)
);
fnc_RTD2456 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100110011000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2456)
);
fnc_RTD2457 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100110011001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2457)
);
fnc_RTD2458 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100110011010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2458)
);
fnc_RTD2459 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100110011011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2459)
);
fnc_RTD2460 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100110011100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2460)
);
fnc_RTD2461 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100110011101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2461)
);
fnc_RTD2462 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100110011110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2462)
);
fnc_RTD2463 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100110011111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2463)
);
fnc_RTD2464 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100110100000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2464)
);
fnc_RTD2465 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100110100001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2465)
);
fnc_RTD2466 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100110100010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2466)
);
fnc_RTD2467 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100110100011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2467)
);
fnc_RTD2468 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100110100100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2468)
);
fnc_RTD2469 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100110100101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2469)
);
fnc_RTD2470 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100110100110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2470)
);
fnc_RTD2471 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100110100111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2471)
);
fnc_RTD2472 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100110101000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2472)
);
fnc_RTD2473 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100110101001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2473)
);
fnc_RTD2474 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100110101010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2474)
);
fnc_RTD2475 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100110101011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2475)
);
fnc_RTD2476 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100110101100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2476)
);
fnc_RTD2477 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100110101101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2477)
);
fnc_RTD2478 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100110101110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2478)
);
fnc_RTD2479 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100110101111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2479)
);
fnc_RTD2480 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100110110000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2480)
);
fnc_RTD2481 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100110110001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2481)
);
fnc_RTD2482 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100110110010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2482)
);
fnc_RTD2483 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100110110011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2483)
);
fnc_RTD2484 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100110110100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2484)
);
fnc_RTD2485 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100110110101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2485)
);
fnc_RTD2486 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100110110110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2486)
);
fnc_RTD2487 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100110110111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2487)
);
fnc_RTD2488 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100110111000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2488)
);
fnc_RTD2489 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100110111001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2489)
);
fnc_RTD2490 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100110111010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2490)
);
fnc_RTD2491 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100110111011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2491)
);
fnc_RTD2492 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100110111100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2492)
);
fnc_RTD2493 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100110111101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2493)
);
fnc_RTD2494 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100110111110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2494)
);
fnc_RTD2495 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100110111111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2495)
);
fnc_RTD2496 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100111000000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2496)
);
fnc_RTD2497 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100111000001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2497)
);
fnc_RTD2498 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100111000010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2498)
);
fnc_RTD2499 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100111000011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2499)
);
fnc_RTD2500 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100111000100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2500)
);
fnc_RTD2501 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100111000101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2501)
);
fnc_RTD2502 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100111000110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2502)
);
fnc_RTD2503 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100111000111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2503)
);
fnc_RTD2504 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100111001000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2504)
);
fnc_RTD2505 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100111001001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2505)
);
fnc_RTD2506 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100111001010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2506)
);
fnc_RTD2507 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100111001011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2507)
);
fnc_RTD2508 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100111001100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2508)
);
fnc_RTD2509 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100111001101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2509)
);
fnc_RTD2510 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100111001110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2510)
);
fnc_RTD2511 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100111001111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2511)
);
fnc_RTD2512 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100111010000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2512)
);
fnc_RTD2513 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100111010001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2513)
);
fnc_RTD2514 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100111010010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2514)
);
fnc_RTD2515 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100111010011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2515)
);
fnc_RTD2516 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100111010100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2516)
);
fnc_RTD2517 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100111010101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2517)
);
fnc_RTD2518 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100111010110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2518)
);
fnc_RTD2519 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100111010111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2519)
);
fnc_RTD2520 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100111011000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2520)
);
fnc_RTD2521 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100111011001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2521)
);
fnc_RTD2522 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100111011010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2522)
);
fnc_RTD2523 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100111011011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2523)
);
fnc_RTD2524 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100111011100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2524)
);
fnc_RTD2525 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100111011101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2525)
);
fnc_RTD2526 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100111011110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2526)
);
fnc_RTD2527 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100111011111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2527)
);
fnc_RTD2528 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100111100000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2528)
);
fnc_RTD2529 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100111100001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2529)
);
fnc_RTD2530 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100111100010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2530)
);
fnc_RTD2531 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100111100011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2531)
);
fnc_RTD2532 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100111100100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2532)
);
fnc_RTD2533 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100111100101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2533)
);
fnc_RTD2534 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100111100110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2534)
);
fnc_RTD2535 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100111100111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2535)
);
fnc_RTD2536 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100111101000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2536)
);
fnc_RTD2537 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100111101001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2537)
);
fnc_RTD2538 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100111101010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2538)
);
fnc_RTD2539 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100111101011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2539)
);
fnc_RTD2540 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100111101100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2540)
);
fnc_RTD2541 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100111101101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2541)
);
fnc_RTD2542 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100111101110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2542)
);
fnc_RTD2543 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100111101111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2543)
);
fnc_RTD2544 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100111110000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2544)
);
fnc_RTD2545 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100111110001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2545)
);
fnc_RTD2546 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100111110010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2546)
);
fnc_RTD2547 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100111110011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2547)
);
fnc_RTD2548 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100111110100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2548)
);
fnc_RTD2549 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100111110101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2549)
);
fnc_RTD2550 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100111110110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2550)
);
fnc_RTD2551 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100111110111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2551)
);
fnc_RTD2552 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100111111000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2552)
);
fnc_RTD2553 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100111111001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2553)
);
fnc_RTD2554 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100111111010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2554)
);
fnc_RTD2555 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100111111011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2555)
);
fnc_RTD2556 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100111111100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2556)
);
fnc_RTD2557 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100111111101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2557)
);
fnc_RTD2558 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100111111110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2558)
);
fnc_RTD2559 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000100111111111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2559)
);
fnc_RTD2560 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101000000000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2560)
);
fnc_RTD2561 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101000000001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2561)
);
fnc_RTD2562 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101000000010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2562)
);
fnc_RTD2563 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101000000011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2563)
);
fnc_RTD2564 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101000000100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2564)
);
fnc_RTD2565 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101000000101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2565)
);
fnc_RTD2566 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101000000110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2566)
);
fnc_RTD2567 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101000000111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2567)
);
fnc_RTD2568 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101000001000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2568)
);
fnc_RTD2569 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101000001001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2569)
);
fnc_RTD2570 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101000001010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2570)
);
fnc_RTD2571 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101000001011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2571)
);
fnc_RTD2572 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101000001100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2572)
);
fnc_RTD2573 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101000001101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2573)
);
fnc_RTD2574 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101000001110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2574)
);
fnc_RTD2575 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101000001111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2575)
);
fnc_RTD2576 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101000010000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2576)
);
fnc_RTD2577 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101000010001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2577)
);
fnc_RTD2578 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101000010010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2578)
);
fnc_RTD2579 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101000010011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2579)
);
fnc_RTD2580 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101000010100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2580)
);
fnc_RTD2581 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101000010101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2581)
);
fnc_RTD2582 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101000010110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2582)
);
fnc_RTD2583 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101000010111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2583)
);
fnc_RTD2584 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101000011000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2584)
);
fnc_RTD2585 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101000011001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2585)
);
fnc_RTD2586 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101000011010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2586)
);
fnc_RTD2587 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101000011011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2587)
);
fnc_RTD2588 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101000011100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2588)
);
fnc_RTD2589 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101000011101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2589)
);
fnc_RTD2590 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101000011110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2590)
);
fnc_RTD2591 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101000011111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2591)
);
fnc_RTD2592 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101000100000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2592)
);
fnc_RTD2593 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101000100001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2593)
);
fnc_RTD2594 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101000100010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2594)
);
fnc_RTD2595 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101000100011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2595)
);
fnc_RTD2596 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101000100100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2596)
);
fnc_RTD2597 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101000100101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2597)
);
fnc_RTD2598 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101000100110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2598)
);
fnc_RTD2599 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101000100111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2599)
);
fnc_RTD2600 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101000101000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2600)
);
fnc_RTD2601 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101000101001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2601)
);
fnc_RTD2602 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101000101010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2602)
);
fnc_RTD2603 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101000101011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2603)
);
fnc_RTD2604 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101000101100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2604)
);
fnc_RTD2605 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101000101101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2605)
);
fnc_RTD2606 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101000101110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2606)
);
fnc_RTD2607 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101000101111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2607)
);
fnc_RTD2608 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101000110000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2608)
);
fnc_RTD2609 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101000110001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2609)
);
fnc_RTD2610 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101000110010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2610)
);
fnc_RTD2611 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101000110011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2611)
);
fnc_RTD2612 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101000110100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2612)
);
fnc_RTD2613 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101000110101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2613)
);
fnc_RTD2614 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101000110110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2614)
);
fnc_RTD2615 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101000110111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2615)
);
fnc_RTD2616 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101000111000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2616)
);
fnc_RTD2617 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101000111001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2617)
);
fnc_RTD2618 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101000111010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2618)
);
fnc_RTD2619 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101000111011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2619)
);
fnc_RTD2620 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101000111100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2620)
);
fnc_RTD2621 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101000111101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2621)
);
fnc_RTD2622 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101000111110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2622)
);
fnc_RTD2623 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101000111111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2623)
);
fnc_RTD2624 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101001000000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2624)
);
fnc_RTD2625 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101001000001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2625)
);
fnc_RTD2626 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101001000010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2626)
);
fnc_RTD2627 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101001000011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2627)
);
fnc_RTD2628 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101001000100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2628)
);
fnc_RTD2629 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101001000101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2629)
);
fnc_RTD2630 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101001000110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2630)
);
fnc_RTD2631 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101001000111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2631)
);
fnc_RTD2632 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101001001000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2632)
);
fnc_RTD2633 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101001001001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2633)
);
fnc_RTD2634 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101001001010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2634)
);
fnc_RTD2635 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101001001011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2635)
);
fnc_RTD2636 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101001001100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2636)
);
fnc_RTD2637 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101001001101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2637)
);
fnc_RTD2638 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101001001110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2638)
);
fnc_RTD2639 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101001001111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2639)
);
fnc_RTD2640 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101001010000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2640)
);
fnc_RTD2641 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101001010001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2641)
);
fnc_RTD2642 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101001010010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2642)
);
fnc_RTD2643 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101001010011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2643)
);
fnc_RTD2644 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101001010100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2644)
);
fnc_RTD2645 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101001010101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2645)
);
fnc_RTD2646 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101001010110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2646)
);
fnc_RTD2647 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101001010111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2647)
);
fnc_RTD2648 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101001011000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2648)
);
fnc_RTD2649 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101001011001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2649)
);
fnc_RTD2650 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101001011010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2650)
);
fnc_RTD2651 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101001011011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2651)
);
fnc_RTD2652 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101001011100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2652)
);
fnc_RTD2653 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101001011101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2653)
);
fnc_RTD2654 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101001011110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2654)
);
fnc_RTD2655 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101001011111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2655)
);
fnc_RTD2656 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101001100000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2656)
);
fnc_RTD2657 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101001100001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2657)
);
fnc_RTD2658 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101001100010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2658)
);
fnc_RTD2659 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101001100011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2659)
);
fnc_RTD2660 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101001100100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2660)
);
fnc_RTD2661 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101001100101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2661)
);
fnc_RTD2662 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101001100110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2662)
);
fnc_RTD2663 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101001100111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2663)
);
fnc_RTD2664 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101001101000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2664)
);
fnc_RTD2665 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101001101001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2665)
);
fnc_RTD2666 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101001101010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2666)
);
fnc_RTD2667 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101001101011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2667)
);
fnc_RTD2668 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101001101100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2668)
);
fnc_RTD2669 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101001101101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2669)
);
fnc_RTD2670 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101001101110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2670)
);
fnc_RTD2671 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101001101111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2671)
);
fnc_RTD2672 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101001110000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2672)
);
fnc_RTD2673 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101001110001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2673)
);
fnc_RTD2674 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101001110010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2674)
);
fnc_RTD2675 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101001110011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2675)
);
fnc_RTD2676 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101001110100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2676)
);
fnc_RTD2677 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101001110101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2677)
);
fnc_RTD2678 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101001110110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2678)
);
fnc_RTD2679 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101001110111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2679)
);
fnc_RTD2680 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101001111000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2680)
);
fnc_RTD2681 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101001111001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2681)
);
fnc_RTD2682 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101001111010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2682)
);
fnc_RTD2683 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101001111011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2683)
);
fnc_RTD2684 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101001111100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2684)
);
fnc_RTD2685 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101001111101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2685)
);
fnc_RTD2686 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101001111110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2686)
);
fnc_RTD2687 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101001111111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2687)
);
fnc_RTD2688 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101010000000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2688)
);
fnc_RTD2689 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101010000001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2689)
);
fnc_RTD2690 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101010000010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2690)
);
fnc_RTD2691 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101010000011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2691)
);
fnc_RTD2692 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101010000100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2692)
);
fnc_RTD2693 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101010000101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2693)
);
fnc_RTD2694 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101010000110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2694)
);
fnc_RTD2695 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101010000111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2695)
);
fnc_RTD2696 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101010001000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2696)
);
fnc_RTD2697 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101010001001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2697)
);
fnc_RTD2698 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101010001010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2698)
);
fnc_RTD2699 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101010001011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2699)
);
fnc_RTD2700 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101010001100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2700)
);
fnc_RTD2701 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101010001101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2701)
);
fnc_RTD2702 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101010001110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2702)
);
fnc_RTD2703 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101010001111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2703)
);
fnc_RTD2704 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101010010000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2704)
);
fnc_RTD2705 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101010010001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2705)
);
fnc_RTD2706 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101010010010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2706)
);
fnc_RTD2707 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101010010011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2707)
);
fnc_RTD2708 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101010010100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2708)
);
fnc_RTD2709 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101010010101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2709)
);
fnc_RTD2710 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101010010110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2710)
);
fnc_RTD2711 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101010010111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2711)
);
fnc_RTD2712 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101010011000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2712)
);
fnc_RTD2713 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101010011001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2713)
);
fnc_RTD2714 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101010011010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2714)
);
fnc_RTD2715 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101010011011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2715)
);
fnc_RTD2716 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101010011100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2716)
);
fnc_RTD2717 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101010011101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2717)
);
fnc_RTD2718 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101010011110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2718)
);
fnc_RTD2719 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101010011111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2719)
);
fnc_RTD2720 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101010100000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2720)
);
fnc_RTD2721 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101010100001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2721)
);
fnc_RTD2722 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101010100010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2722)
);
fnc_RTD2723 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101010100011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2723)
);
fnc_RTD2724 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101010100100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2724)
);
fnc_RTD2725 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101010100101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2725)
);
fnc_RTD2726 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101010100110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2726)
);
fnc_RTD2727 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101010100111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2727)
);
fnc_RTD2728 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101010101000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2728)
);
fnc_RTD2729 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101010101001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2729)
);
fnc_RTD2730 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101010101010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2730)
);
fnc_RTD2731 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101010101011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2731)
);
fnc_RTD2732 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101010101100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2732)
);
fnc_RTD2733 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101010101101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2733)
);
fnc_RTD2734 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101010101110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2734)
);
fnc_RTD2735 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101010101111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2735)
);
fnc_RTD2736 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101010110000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2736)
);
fnc_RTD2737 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101010110001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2737)
);
fnc_RTD2738 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101010110010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2738)
);
fnc_RTD2739 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101010110011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2739)
);
fnc_RTD2740 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101010110100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2740)
);
fnc_RTD2741 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101010110101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2741)
);
fnc_RTD2742 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101010110110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2742)
);
fnc_RTD2743 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101010110111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2743)
);
fnc_RTD2744 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101010111000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2744)
);
fnc_RTD2745 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101010111001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2745)
);
fnc_RTD2746 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101010111010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2746)
);
fnc_RTD2747 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101010111011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2747)
);
fnc_RTD2748 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101010111100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2748)
);
fnc_RTD2749 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101010111101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2749)
);
fnc_RTD2750 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101010111110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2750)
);
fnc_RTD2751 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101010111111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2751)
);
fnc_RTD2752 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101011000000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2752)
);
fnc_RTD2753 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101011000001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2753)
);
fnc_RTD2754 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101011000010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2754)
);
fnc_RTD2755 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101011000011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2755)
);
fnc_RTD2756 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101011000100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2756)
);
fnc_RTD2757 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101011000101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2757)
);
fnc_RTD2758 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101011000110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2758)
);
fnc_RTD2759 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101011000111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2759)
);
fnc_RTD2760 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101011001000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2760)
);
fnc_RTD2761 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101011001001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2761)
);
fnc_RTD2762 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101011001010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2762)
);
fnc_RTD2763 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101011001011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2763)
);
fnc_RTD2764 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101011001100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2764)
);
fnc_RTD2765 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101011001101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2765)
);
fnc_RTD2766 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101011001110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2766)
);
fnc_RTD2767 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101011001111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2767)
);
fnc_RTD2768 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101011010000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2768)
);
fnc_RTD2769 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101011010001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2769)
);
fnc_RTD2770 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101011010010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2770)
);
fnc_RTD2771 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101011010011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2771)
);
fnc_RTD2772 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101011010100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2772)
);
fnc_RTD2773 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101011010101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2773)
);
fnc_RTD2774 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101011010110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2774)
);
fnc_RTD2775 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101011010111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2775)
);
fnc_RTD2776 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101011011000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2776)
);
fnc_RTD2777 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101011011001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2777)
);
fnc_RTD2778 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101011011010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2778)
);
fnc_RTD2779 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101011011011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2779)
);
fnc_RTD2780 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101011011100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2780)
);
fnc_RTD2781 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101011011101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2781)
);
fnc_RTD2782 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101011011110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2782)
);
fnc_RTD2783 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101011011111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2783)
);
fnc_RTD2784 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101011100000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2784)
);
fnc_RTD2785 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101011100001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2785)
);
fnc_RTD2786 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101011100010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2786)
);
fnc_RTD2787 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101011100011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2787)
);
fnc_RTD2788 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101011100100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2788)
);
fnc_RTD2789 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101011100101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2789)
);
fnc_RTD2790 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101011100110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2790)
);
fnc_RTD2791 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101011100111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2791)
);
fnc_RTD2792 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101011101000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2792)
);
fnc_RTD2793 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101011101001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2793)
);
fnc_RTD2794 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101011101010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2794)
);
fnc_RTD2795 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101011101011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2795)
);
fnc_RTD2796 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101011101100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2796)
);
fnc_RTD2797 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101011101101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2797)
);
fnc_RTD2798 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101011101110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2798)
);
fnc_RTD2799 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000101011101111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_RTD),
	match_result_o      => sig_fnc_RTD(2799)
);
bram_VERS : xilinx_single_port_ram_no_change generic map (
	RAM_WIDTH => C_BRAM_VERS_WIDTH,
	RAM_DEPTH => C_BRAM_VERS_DEPTH,
	RAM_PERFORMANCE => "LOW_LATENCY", --"HIGH_PERFORMANCE",
	INIT_FILE => "bram_VERS.mem"
) port map (
	clka   => clk_i,
	addra  => query_i(C_QUERY_VERS)((clogb2(C_BRAM_VERS_DEPTH)-1) downto 0),
	dina   => mem_i(C_BRAM_VERS_WIDTH-1 downto 0),
	wea    => meme_i(C_BRAM_VERS),
	ena    => '1',
	rsta   => '0',
	regcea => '1',
	douta  => sig_ram_VERS
);
fnc_OWN0 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000000000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(0)
);
fnc_OWN1 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000000001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1)
);
fnc_OWN2 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000000010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(2)
);
fnc_OWN3 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000000011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(3)
);
fnc_OWN4 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000000100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(4)
);
fnc_OWN5 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000000101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(5)
);
fnc_OWN6 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000000110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(6)
);
fnc_OWN7 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000000111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(7)
);
fnc_OWN8 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000001000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(8)
);
fnc_OWN9 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000001001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(9)
);
fnc_OWN10 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000001010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(10)
);
fnc_OWN11 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000001011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(11)
);
fnc_OWN12 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000001100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(12)
);
fnc_OWN13 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000001101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(13)
);
fnc_OWN14 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000001110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(14)
);
fnc_OWN15 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000001111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(15)
);
fnc_OWN16 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000010000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(16)
);
fnc_OWN17 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000010001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(17)
);
fnc_OWN18 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000010010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(18)
);
fnc_OWN19 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000010011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(19)
);
fnc_OWN20 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000010100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(20)
);
fnc_OWN21 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000010101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(21)
);
fnc_OWN22 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000010110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(22)
);
fnc_OWN23 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000010111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(23)
);
fnc_OWN24 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000011000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(24)
);
fnc_OWN25 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000011001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(25)
);
fnc_OWN26 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000011010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(26)
);
fnc_OWN27 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000011011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(27)
);
fnc_OWN28 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000011100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(28)
);
fnc_OWN29 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000011101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(29)
);
fnc_OWN30 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000011110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(30)
);
fnc_OWN31 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000011111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(31)
);
fnc_OWN32 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000100000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(32)
);
fnc_OWN33 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000100001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(33)
);
fnc_OWN34 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000100010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(34)
);
fnc_OWN35 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000100011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(35)
);
fnc_OWN36 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000100100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(36)
);
fnc_OWN37 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000100101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(37)
);
fnc_OWN38 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000100110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(38)
);
fnc_OWN39 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000100111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(39)
);
fnc_OWN40 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000101000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(40)
);
fnc_OWN41 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000101001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(41)
);
fnc_OWN42 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000101010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(42)
);
fnc_OWN43 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000101011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(43)
);
fnc_OWN44 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000101100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(44)
);
fnc_OWN45 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000101101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(45)
);
fnc_OWN46 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000101110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(46)
);
fnc_OWN47 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000101111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(47)
);
fnc_OWN48 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000110000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(48)
);
fnc_OWN49 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000110001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(49)
);
fnc_OWN50 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000110010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(50)
);
fnc_OWN51 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000110011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(51)
);
fnc_OWN52 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000110100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(52)
);
fnc_OWN53 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000110101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(53)
);
fnc_OWN54 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000110110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(54)
);
fnc_OWN55 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000110111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(55)
);
fnc_OWN56 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000111000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(56)
);
fnc_OWN57 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000111001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(57)
);
fnc_OWN58 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000111010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(58)
);
fnc_OWN59 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000111011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(59)
);
fnc_OWN60 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000111100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(60)
);
fnc_OWN61 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000111101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(61)
);
fnc_OWN62 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000111110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(62)
);
fnc_OWN63 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000000111111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(63)
);
fnc_OWN64 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001000000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(64)
);
fnc_OWN65 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001000001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(65)
);
fnc_OWN66 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001000010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(66)
);
fnc_OWN67 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001000011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(67)
);
fnc_OWN68 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001000100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(68)
);
fnc_OWN69 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001000101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(69)
);
fnc_OWN70 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001000110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(70)
);
fnc_OWN71 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001000111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(71)
);
fnc_OWN72 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001001000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(72)
);
fnc_OWN73 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001001001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(73)
);
fnc_OWN74 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001001010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(74)
);
fnc_OWN75 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001001011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(75)
);
fnc_OWN76 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001001100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(76)
);
fnc_OWN77 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001001101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(77)
);
fnc_OWN78 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001001110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(78)
);
fnc_OWN79 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001001111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(79)
);
fnc_OWN80 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001010000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(80)
);
fnc_OWN81 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001010001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(81)
);
fnc_OWN82 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001010010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(82)
);
fnc_OWN83 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001010011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(83)
);
fnc_OWN84 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001010100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(84)
);
fnc_OWN85 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001010101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(85)
);
fnc_OWN86 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001010110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(86)
);
fnc_OWN87 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001010111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(87)
);
fnc_OWN88 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001011000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(88)
);
fnc_OWN89 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001011001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(89)
);
fnc_OWN90 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001011010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(90)
);
fnc_OWN91 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001011011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(91)
);
fnc_OWN92 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001011100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(92)
);
fnc_OWN93 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001011101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(93)
);
fnc_OWN94 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001011110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(94)
);
fnc_OWN95 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001011111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(95)
);
fnc_OWN96 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001100000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(96)
);
fnc_OWN97 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001100001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(97)
);
fnc_OWN98 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001100010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(98)
);
fnc_OWN99 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001100011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(99)
);
fnc_OWN100 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001100100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(100)
);
fnc_OWN101 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001100101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(101)
);
fnc_OWN102 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001100110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(102)
);
fnc_OWN103 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001100111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(103)
);
fnc_OWN104 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001101000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(104)
);
fnc_OWN105 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001101001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(105)
);
fnc_OWN106 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001101010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(106)
);
fnc_OWN107 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001101011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(107)
);
fnc_OWN108 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001101100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(108)
);
fnc_OWN109 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001101101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(109)
);
fnc_OWN110 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001101110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(110)
);
fnc_OWN111 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001101111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(111)
);
fnc_OWN112 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001110000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(112)
);
fnc_OWN113 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001110001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(113)
);
fnc_OWN114 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001110010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(114)
);
fnc_OWN115 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001110011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(115)
);
fnc_OWN116 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001110100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(116)
);
fnc_OWN117 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001110101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(117)
);
fnc_OWN118 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001110110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(118)
);
fnc_OWN119 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001110111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(119)
);
fnc_OWN120 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001111000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(120)
);
fnc_OWN121 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001111001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(121)
);
fnc_OWN122 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001111010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(122)
);
fnc_OWN123 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001111011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(123)
);
fnc_OWN124 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001111100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(124)
);
fnc_OWN125 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001111101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(125)
);
fnc_OWN126 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001111110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(126)
);
fnc_OWN127 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000001111111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(127)
);
fnc_OWN128 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010000000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(128)
);
fnc_OWN129 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010000001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(129)
);
fnc_OWN130 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010000010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(130)
);
fnc_OWN131 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010000011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(131)
);
fnc_OWN132 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010000100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(132)
);
fnc_OWN133 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010000101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(133)
);
fnc_OWN134 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010000110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(134)
);
fnc_OWN135 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010000111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(135)
);
fnc_OWN136 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010001000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(136)
);
fnc_OWN137 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010001001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(137)
);
fnc_OWN138 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010001010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(138)
);
fnc_OWN139 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010001011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(139)
);
fnc_OWN140 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010001100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(140)
);
fnc_OWN141 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010001101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(141)
);
fnc_OWN142 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010001110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(142)
);
fnc_OWN143 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010001111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(143)
);
fnc_OWN144 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010010000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(144)
);
fnc_OWN145 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010010001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(145)
);
fnc_OWN146 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010010010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(146)
);
fnc_OWN147 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010010011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(147)
);
fnc_OWN148 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010010100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(148)
);
fnc_OWN149 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010010101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(149)
);
fnc_OWN150 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010010110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(150)
);
fnc_OWN151 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010010111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(151)
);
fnc_OWN152 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010011000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(152)
);
fnc_OWN153 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010011001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(153)
);
fnc_OWN154 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010011010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(154)
);
fnc_OWN155 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010011011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(155)
);
fnc_OWN156 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010011100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(156)
);
fnc_OWN157 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010011101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(157)
);
fnc_OWN158 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010011110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(158)
);
fnc_OWN159 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010011111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(159)
);
fnc_OWN160 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010100000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(160)
);
fnc_OWN161 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010100001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(161)
);
fnc_OWN162 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010100010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(162)
);
fnc_OWN163 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010100011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(163)
);
fnc_OWN164 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010100100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(164)
);
fnc_OWN165 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010100101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(165)
);
fnc_OWN166 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010100110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(166)
);
fnc_OWN167 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010100111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(167)
);
fnc_OWN168 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010101000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(168)
);
fnc_OWN169 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010101001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(169)
);
fnc_OWN170 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010101010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(170)
);
fnc_OWN171 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010101011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(171)
);
fnc_OWN172 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010101100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(172)
);
fnc_OWN173 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010101101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(173)
);
fnc_OWN174 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010101110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(174)
);
fnc_OWN175 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010101111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(175)
);
fnc_OWN176 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010110000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(176)
);
fnc_OWN177 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010110001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(177)
);
fnc_OWN178 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010110010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(178)
);
fnc_OWN179 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010110011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(179)
);
fnc_OWN180 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010110100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(180)
);
fnc_OWN181 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010110101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(181)
);
fnc_OWN182 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010110110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(182)
);
fnc_OWN183 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010110111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(183)
);
fnc_OWN184 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010111000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(184)
);
fnc_OWN185 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010111001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(185)
);
fnc_OWN186 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010111010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(186)
);
fnc_OWN187 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010111011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(187)
);
fnc_OWN188 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010111100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(188)
);
fnc_OWN189 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010111101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(189)
);
fnc_OWN190 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010111110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(190)
);
fnc_OWN191 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000010111111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(191)
);
fnc_OWN192 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011000000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(192)
);
fnc_OWN193 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011000001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(193)
);
fnc_OWN194 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011000010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(194)
);
fnc_OWN195 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011000011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(195)
);
fnc_OWN196 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011000100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(196)
);
fnc_OWN197 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011000101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(197)
);
fnc_OWN198 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011000110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(198)
);
fnc_OWN199 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011000111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(199)
);
fnc_OWN200 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011001000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(200)
);
fnc_OWN201 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011001001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(201)
);
fnc_OWN202 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011001010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(202)
);
fnc_OWN203 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011001011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(203)
);
fnc_OWN204 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011001100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(204)
);
fnc_OWN205 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011001101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(205)
);
fnc_OWN206 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011001110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(206)
);
fnc_OWN207 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011001111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(207)
);
fnc_OWN208 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011010000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(208)
);
fnc_OWN209 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011010001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(209)
);
fnc_OWN210 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011010010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(210)
);
fnc_OWN211 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011010011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(211)
);
fnc_OWN212 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011010100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(212)
);
fnc_OWN213 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011010101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(213)
);
fnc_OWN214 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011010110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(214)
);
fnc_OWN215 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011010111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(215)
);
fnc_OWN216 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011011000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(216)
);
fnc_OWN217 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011011001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(217)
);
fnc_OWN218 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011011010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(218)
);
fnc_OWN219 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011011011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(219)
);
fnc_OWN220 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011011100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(220)
);
fnc_OWN221 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011011101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(221)
);
fnc_OWN222 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011011110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(222)
);
fnc_OWN223 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011011111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(223)
);
fnc_OWN224 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011100000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(224)
);
fnc_OWN225 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011100001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(225)
);
fnc_OWN226 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011100010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(226)
);
fnc_OWN227 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011100011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(227)
);
fnc_OWN228 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011100100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(228)
);
fnc_OWN229 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011100101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(229)
);
fnc_OWN230 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011100110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(230)
);
fnc_OWN231 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011100111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(231)
);
fnc_OWN232 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011101000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(232)
);
fnc_OWN233 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011101001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(233)
);
fnc_OWN234 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011101010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(234)
);
fnc_OWN235 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011101011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(235)
);
fnc_OWN236 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011101100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(236)
);
fnc_OWN237 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011101101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(237)
);
fnc_OWN238 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011101110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(238)
);
fnc_OWN239 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011101111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(239)
);
fnc_OWN240 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011110000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(240)
);
fnc_OWN241 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011110001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(241)
);
fnc_OWN242 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011110010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(242)
);
fnc_OWN243 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011110011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(243)
);
fnc_OWN244 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011110100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(244)
);
fnc_OWN245 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011110101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(245)
);
fnc_OWN246 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011110110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(246)
);
fnc_OWN247 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011110111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(247)
);
fnc_OWN248 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011111000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(248)
);
fnc_OWN249 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011111001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(249)
);
fnc_OWN250 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011111010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(250)
);
fnc_OWN251 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011111011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(251)
);
fnc_OWN252 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011111100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(252)
);
fnc_OWN253 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011111101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(253)
);
fnc_OWN254 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011111110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(254)
);
fnc_OWN255 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000011111111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(255)
);
fnc_OWN256 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100000000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(256)
);
fnc_OWN257 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100000001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(257)
);
fnc_OWN258 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100000010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(258)
);
fnc_OWN259 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100000011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(259)
);
fnc_OWN260 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100000100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(260)
);
fnc_OWN261 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100000101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(261)
);
fnc_OWN262 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100000110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(262)
);
fnc_OWN263 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100000111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(263)
);
fnc_OWN264 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100001000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(264)
);
fnc_OWN265 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100001001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(265)
);
fnc_OWN266 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100001010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(266)
);
fnc_OWN267 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100001011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(267)
);
fnc_OWN268 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100001100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(268)
);
fnc_OWN269 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100001101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(269)
);
fnc_OWN270 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100001110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(270)
);
fnc_OWN271 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100001111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(271)
);
fnc_OWN272 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100010000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(272)
);
fnc_OWN273 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100010001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(273)
);
fnc_OWN274 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100010010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(274)
);
fnc_OWN275 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100010011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(275)
);
fnc_OWN276 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100010100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(276)
);
fnc_OWN277 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100010101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(277)
);
fnc_OWN278 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100010110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(278)
);
fnc_OWN279 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100010111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(279)
);
fnc_OWN280 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100011000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(280)
);
fnc_OWN281 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100011001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(281)
);
fnc_OWN282 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100011010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(282)
);
fnc_OWN283 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100011011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(283)
);
fnc_OWN284 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100011100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(284)
);
fnc_OWN285 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100011101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(285)
);
fnc_OWN286 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100011110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(286)
);
fnc_OWN287 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100011111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(287)
);
fnc_OWN288 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100100000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(288)
);
fnc_OWN289 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100100001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(289)
);
fnc_OWN290 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100100010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(290)
);
fnc_OWN291 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100100011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(291)
);
fnc_OWN292 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100100100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(292)
);
fnc_OWN293 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100100101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(293)
);
fnc_OWN294 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100100110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(294)
);
fnc_OWN295 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100100111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(295)
);
fnc_OWN296 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100101000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(296)
);
fnc_OWN297 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100101001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(297)
);
fnc_OWN298 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100101010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(298)
);
fnc_OWN299 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100101011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(299)
);
fnc_OWN300 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100101100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(300)
);
fnc_OWN301 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100101101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(301)
);
fnc_OWN302 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100101110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(302)
);
fnc_OWN303 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100101111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(303)
);
fnc_OWN304 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100110000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(304)
);
fnc_OWN305 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100110001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(305)
);
fnc_OWN306 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100110010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(306)
);
fnc_OWN307 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100110011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(307)
);
fnc_OWN308 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100110100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(308)
);
fnc_OWN309 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100110101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(309)
);
fnc_OWN310 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100110110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(310)
);
fnc_OWN311 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100110111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(311)
);
fnc_OWN312 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100111000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(312)
);
fnc_OWN313 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100111001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(313)
);
fnc_OWN314 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100111010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(314)
);
fnc_OWN315 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100111011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(315)
);
fnc_OWN316 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100111100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(316)
);
fnc_OWN317 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100111101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(317)
);
fnc_OWN318 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100111110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(318)
);
fnc_OWN319 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000100111111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(319)
);
fnc_OWN320 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101000000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(320)
);
fnc_OWN321 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101000001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(321)
);
fnc_OWN322 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101000010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(322)
);
fnc_OWN323 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101000011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(323)
);
fnc_OWN324 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101000100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(324)
);
fnc_OWN325 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101000101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(325)
);
fnc_OWN326 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101000110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(326)
);
fnc_OWN327 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101000111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(327)
);
fnc_OWN328 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101001000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(328)
);
fnc_OWN329 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101001001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(329)
);
fnc_OWN330 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101001010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(330)
);
fnc_OWN331 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101001011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(331)
);
fnc_OWN332 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101001100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(332)
);
fnc_OWN333 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101001101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(333)
);
fnc_OWN334 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101001110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(334)
);
fnc_OWN335 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101001111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(335)
);
fnc_OWN336 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101010000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(336)
);
fnc_OWN337 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101010001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(337)
);
fnc_OWN338 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101010010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(338)
);
fnc_OWN339 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101010011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(339)
);
fnc_OWN340 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101010100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(340)
);
fnc_OWN341 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101010101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(341)
);
fnc_OWN342 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101010110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(342)
);
fnc_OWN343 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101010111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(343)
);
fnc_OWN344 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101011000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(344)
);
fnc_OWN345 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101011001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(345)
);
fnc_OWN346 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101011010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(346)
);
fnc_OWN347 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101011011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(347)
);
fnc_OWN348 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101011100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(348)
);
fnc_OWN349 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101011101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(349)
);
fnc_OWN350 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101011110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(350)
);
fnc_OWN351 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101011111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(351)
);
fnc_OWN352 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101100000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(352)
);
fnc_OWN353 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101100001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(353)
);
fnc_OWN354 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101100010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(354)
);
fnc_OWN355 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101100011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(355)
);
fnc_OWN356 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101100100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(356)
);
fnc_OWN357 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101100101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(357)
);
fnc_OWN358 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101100110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(358)
);
fnc_OWN359 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101100111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(359)
);
fnc_OWN360 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101101000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(360)
);
fnc_OWN361 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101101001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(361)
);
fnc_OWN362 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101101010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(362)
);
fnc_OWN363 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101101011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(363)
);
fnc_OWN364 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101101100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(364)
);
fnc_OWN365 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101101101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(365)
);
fnc_OWN366 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101101110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(366)
);
fnc_OWN367 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101101111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(367)
);
fnc_OWN368 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101110000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(368)
);
fnc_OWN369 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101110001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(369)
);
fnc_OWN370 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101110010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(370)
);
fnc_OWN371 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101110011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(371)
);
fnc_OWN372 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101110100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(372)
);
fnc_OWN373 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101110101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(373)
);
fnc_OWN374 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101110110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(374)
);
fnc_OWN375 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101110111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(375)
);
fnc_OWN376 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101111000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(376)
);
fnc_OWN377 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101111001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(377)
);
fnc_OWN378 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101111010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(378)
);
fnc_OWN379 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101111011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(379)
);
fnc_OWN380 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101111100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(380)
);
fnc_OWN381 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101111101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(381)
);
fnc_OWN382 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101111110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(382)
);
fnc_OWN383 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000101111111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(383)
);
fnc_OWN384 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110000000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(384)
);
fnc_OWN385 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110000001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(385)
);
fnc_OWN386 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110000010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(386)
);
fnc_OWN387 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110000011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(387)
);
fnc_OWN388 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110000100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(388)
);
fnc_OWN389 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110000101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(389)
);
fnc_OWN390 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110000110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(390)
);
fnc_OWN391 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110000111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(391)
);
fnc_OWN392 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110001000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(392)
);
fnc_OWN393 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110001001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(393)
);
fnc_OWN394 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110001010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(394)
);
fnc_OWN395 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110001011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(395)
);
fnc_OWN396 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110001100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(396)
);
fnc_OWN397 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110001101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(397)
);
fnc_OWN398 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110001110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(398)
);
fnc_OWN399 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110001111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(399)
);
fnc_OWN400 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110010000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(400)
);
fnc_OWN401 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110010001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(401)
);
fnc_OWN402 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110010010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(402)
);
fnc_OWN403 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110010011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(403)
);
fnc_OWN404 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110010100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(404)
);
fnc_OWN405 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110010101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(405)
);
fnc_OWN406 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110010110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(406)
);
fnc_OWN407 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110010111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(407)
);
fnc_OWN408 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110011000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(408)
);
fnc_OWN409 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110011001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(409)
);
fnc_OWN410 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110011010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(410)
);
fnc_OWN411 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110011011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(411)
);
fnc_OWN412 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110011100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(412)
);
fnc_OWN413 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110011101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(413)
);
fnc_OWN414 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110011110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(414)
);
fnc_OWN415 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110011111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(415)
);
fnc_OWN416 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110100000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(416)
);
fnc_OWN417 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110100001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(417)
);
fnc_OWN418 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110100010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(418)
);
fnc_OWN419 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110100011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(419)
);
fnc_OWN420 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110100100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(420)
);
fnc_OWN421 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110100101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(421)
);
fnc_OWN422 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110100110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(422)
);
fnc_OWN423 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110100111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(423)
);
fnc_OWN424 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110101000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(424)
);
fnc_OWN425 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110101001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(425)
);
fnc_OWN426 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110101010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(426)
);
fnc_OWN427 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110101011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(427)
);
fnc_OWN428 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110101100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(428)
);
fnc_OWN429 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110101101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(429)
);
fnc_OWN430 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110101110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(430)
);
fnc_OWN431 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110101111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(431)
);
fnc_OWN432 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110110000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(432)
);
fnc_OWN433 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110110001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(433)
);
fnc_OWN434 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110110010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(434)
);
fnc_OWN435 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110110011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(435)
);
fnc_OWN436 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110110100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(436)
);
fnc_OWN437 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110110101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(437)
);
fnc_OWN438 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110110110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(438)
);
fnc_OWN439 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110110111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(439)
);
fnc_OWN440 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110111000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(440)
);
fnc_OWN441 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110111001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(441)
);
fnc_OWN442 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110111010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(442)
);
fnc_OWN443 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110111011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(443)
);
fnc_OWN444 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110111100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(444)
);
fnc_OWN445 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110111101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(445)
);
fnc_OWN446 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110111110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(446)
);
fnc_OWN447 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000110111111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(447)
);
fnc_OWN448 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111000000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(448)
);
fnc_OWN449 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111000001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(449)
);
fnc_OWN450 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111000010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(450)
);
fnc_OWN451 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111000011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(451)
);
fnc_OWN452 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111000100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(452)
);
fnc_OWN453 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111000101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(453)
);
fnc_OWN454 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111000110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(454)
);
fnc_OWN455 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111000111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(455)
);
fnc_OWN456 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111001000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(456)
);
fnc_OWN457 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111001001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(457)
);
fnc_OWN458 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111001010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(458)
);
fnc_OWN459 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111001011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(459)
);
fnc_OWN460 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111001100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(460)
);
fnc_OWN461 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111001101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(461)
);
fnc_OWN462 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111001110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(462)
);
fnc_OWN463 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111001111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(463)
);
fnc_OWN464 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111010000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(464)
);
fnc_OWN465 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111010001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(465)
);
fnc_OWN466 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111010010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(466)
);
fnc_OWN467 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111010011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(467)
);
fnc_OWN468 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111010100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(468)
);
fnc_OWN469 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111010101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(469)
);
fnc_OWN470 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111010110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(470)
);
fnc_OWN471 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111010111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(471)
);
fnc_OWN472 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111011000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(472)
);
fnc_OWN473 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111011001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(473)
);
fnc_OWN474 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111011010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(474)
);
fnc_OWN475 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111011011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(475)
);
fnc_OWN476 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111011100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(476)
);
fnc_OWN477 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111011101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(477)
);
fnc_OWN478 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111011110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(478)
);
fnc_OWN479 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111011111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(479)
);
fnc_OWN480 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111100000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(480)
);
fnc_OWN481 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111100001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(481)
);
fnc_OWN482 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111100010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(482)
);
fnc_OWN483 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111100011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(483)
);
fnc_OWN484 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111100100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(484)
);
fnc_OWN485 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111100101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(485)
);
fnc_OWN486 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111100110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(486)
);
fnc_OWN487 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111100111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(487)
);
fnc_OWN488 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111101000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(488)
);
fnc_OWN489 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111101001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(489)
);
fnc_OWN490 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111101010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(490)
);
fnc_OWN491 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111101011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(491)
);
fnc_OWN492 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111101100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(492)
);
fnc_OWN493 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111101101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(493)
);
fnc_OWN494 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111101110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(494)
);
fnc_OWN495 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111101111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(495)
);
fnc_OWN496 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111110000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(496)
);
fnc_OWN497 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111110001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(497)
);
fnc_OWN498 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111110010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(498)
);
fnc_OWN499 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111110011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(499)
);
fnc_OWN500 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111110100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(500)
);
fnc_OWN501 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111110101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(501)
);
fnc_OWN502 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111110110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(502)
);
fnc_OWN503 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111110111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(503)
);
fnc_OWN504 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111111000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(504)
);
fnc_OWN505 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111111001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(505)
);
fnc_OWN506 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111111010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(506)
);
fnc_OWN507 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111111011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(507)
);
fnc_OWN508 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111111100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(508)
);
fnc_OWN509 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111111101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(509)
);
fnc_OWN510 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111111110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(510)
);
fnc_OWN511 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000000111111111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(511)
);
fnc_OWN512 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000000000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(512)
);
fnc_OWN513 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000000001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(513)
);
fnc_OWN514 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000000010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(514)
);
fnc_OWN515 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000000011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(515)
);
fnc_OWN516 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000000100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(516)
);
fnc_OWN517 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000000101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(517)
);
fnc_OWN518 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000000110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(518)
);
fnc_OWN519 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000000111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(519)
);
fnc_OWN520 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000001000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(520)
);
fnc_OWN521 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000001001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(521)
);
fnc_OWN522 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000001010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(522)
);
fnc_OWN523 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000001011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(523)
);
fnc_OWN524 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000001100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(524)
);
fnc_OWN525 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000001101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(525)
);
fnc_OWN526 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000001110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(526)
);
fnc_OWN527 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000001111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(527)
);
fnc_OWN528 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000010000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(528)
);
fnc_OWN529 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000010001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(529)
);
fnc_OWN530 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000010010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(530)
);
fnc_OWN531 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000010011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(531)
);
fnc_OWN532 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000010100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(532)
);
fnc_OWN533 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000010101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(533)
);
fnc_OWN534 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000010110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(534)
);
fnc_OWN535 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000010111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(535)
);
fnc_OWN536 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000011000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(536)
);
fnc_OWN537 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000011001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(537)
);
fnc_OWN538 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000011010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(538)
);
fnc_OWN539 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000011011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(539)
);
fnc_OWN540 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000011100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(540)
);
fnc_OWN541 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000011101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(541)
);
fnc_OWN542 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000011110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(542)
);
fnc_OWN543 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000011111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(543)
);
fnc_OWN544 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000100000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(544)
);
fnc_OWN545 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000100001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(545)
);
fnc_OWN546 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000100010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(546)
);
fnc_OWN547 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000100011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(547)
);
fnc_OWN548 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000100100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(548)
);
fnc_OWN549 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000100101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(549)
);
fnc_OWN550 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000100110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(550)
);
fnc_OWN551 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000100111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(551)
);
fnc_OWN552 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000101000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(552)
);
fnc_OWN553 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000101001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(553)
);
fnc_OWN554 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000101010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(554)
);
fnc_OWN555 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000101011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(555)
);
fnc_OWN556 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000101100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(556)
);
fnc_OWN557 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000101101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(557)
);
fnc_OWN558 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000101110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(558)
);
fnc_OWN559 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000101111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(559)
);
fnc_OWN560 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000110000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(560)
);
fnc_OWN561 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000110001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(561)
);
fnc_OWN562 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000110010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(562)
);
fnc_OWN563 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000110011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(563)
);
fnc_OWN564 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000110100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(564)
);
fnc_OWN565 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000110101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(565)
);
fnc_OWN566 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000110110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(566)
);
fnc_OWN567 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000110111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(567)
);
fnc_OWN568 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000111000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(568)
);
fnc_OWN569 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000111001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(569)
);
fnc_OWN570 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000111010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(570)
);
fnc_OWN571 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000111011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(571)
);
fnc_OWN572 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000111100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(572)
);
fnc_OWN573 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000111101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(573)
);
fnc_OWN574 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000111110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(574)
);
fnc_OWN575 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001000111111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(575)
);
fnc_OWN576 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001000000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(576)
);
fnc_OWN577 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001000001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(577)
);
fnc_OWN578 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001000010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(578)
);
fnc_OWN579 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001000011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(579)
);
fnc_OWN580 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001000100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(580)
);
fnc_OWN581 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001000101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(581)
);
fnc_OWN582 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001000110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(582)
);
fnc_OWN583 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001000111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(583)
);
fnc_OWN584 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001001000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(584)
);
fnc_OWN585 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001001001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(585)
);
fnc_OWN586 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001001010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(586)
);
fnc_OWN587 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001001011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(587)
);
fnc_OWN588 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001001100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(588)
);
fnc_OWN589 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001001101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(589)
);
fnc_OWN590 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001001110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(590)
);
fnc_OWN591 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001001111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(591)
);
fnc_OWN592 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001010000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(592)
);
fnc_OWN593 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001010001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(593)
);
fnc_OWN594 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001010010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(594)
);
fnc_OWN595 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001010011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(595)
);
fnc_OWN596 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001010100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(596)
);
fnc_OWN597 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001010101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(597)
);
fnc_OWN598 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001010110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(598)
);
fnc_OWN599 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001010111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(599)
);
fnc_OWN600 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001011000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(600)
);
fnc_OWN601 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001011001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(601)
);
fnc_OWN602 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001011010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(602)
);
fnc_OWN603 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001011011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(603)
);
fnc_OWN604 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001011100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(604)
);
fnc_OWN605 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001011101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(605)
);
fnc_OWN606 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001011110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(606)
);
fnc_OWN607 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001011111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(607)
);
fnc_OWN608 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001100000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(608)
);
fnc_OWN609 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001100001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(609)
);
fnc_OWN610 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001100010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(610)
);
fnc_OWN611 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001100011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(611)
);
fnc_OWN612 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001100100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(612)
);
fnc_OWN613 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001100101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(613)
);
fnc_OWN614 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001100110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(614)
);
fnc_OWN615 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001100111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(615)
);
fnc_OWN616 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001101000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(616)
);
fnc_OWN617 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001101001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(617)
);
fnc_OWN618 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001101010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(618)
);
fnc_OWN619 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001101011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(619)
);
fnc_OWN620 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001101100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(620)
);
fnc_OWN621 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001101101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(621)
);
fnc_OWN622 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001101110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(622)
);
fnc_OWN623 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001101111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(623)
);
fnc_OWN624 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001110000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(624)
);
fnc_OWN625 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001110001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(625)
);
fnc_OWN626 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001110010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(626)
);
fnc_OWN627 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001110011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(627)
);
fnc_OWN628 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001110100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(628)
);
fnc_OWN629 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001110101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(629)
);
fnc_OWN630 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001110110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(630)
);
fnc_OWN631 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001110111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(631)
);
fnc_OWN632 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001111000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(632)
);
fnc_OWN633 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001111001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(633)
);
fnc_OWN634 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001111010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(634)
);
fnc_OWN635 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001111011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(635)
);
fnc_OWN636 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001111100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(636)
);
fnc_OWN637 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001111101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(637)
);
fnc_OWN638 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001111110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(638)
);
fnc_OWN639 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001001111111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(639)
);
fnc_OWN640 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010000000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(640)
);
fnc_OWN641 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010000001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(641)
);
fnc_OWN642 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010000010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(642)
);
fnc_OWN643 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010000011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(643)
);
fnc_OWN644 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010000100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(644)
);
fnc_OWN645 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010000101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(645)
);
fnc_OWN646 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010000110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(646)
);
fnc_OWN647 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010000111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(647)
);
fnc_OWN648 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010001000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(648)
);
fnc_OWN649 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010001001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(649)
);
fnc_OWN650 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010001010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(650)
);
fnc_OWN651 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010001011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(651)
);
fnc_OWN652 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010001100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(652)
);
fnc_OWN653 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010001101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(653)
);
fnc_OWN654 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010001110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(654)
);
fnc_OWN655 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010001111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(655)
);
fnc_OWN656 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010010000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(656)
);
fnc_OWN657 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010010001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(657)
);
fnc_OWN658 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010010010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(658)
);
fnc_OWN659 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010010011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(659)
);
fnc_OWN660 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010010100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(660)
);
fnc_OWN661 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010010101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(661)
);
fnc_OWN662 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010010110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(662)
);
fnc_OWN663 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010010111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(663)
);
fnc_OWN664 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010011000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(664)
);
fnc_OWN665 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010011001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(665)
);
fnc_OWN666 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010011010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(666)
);
fnc_OWN667 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010011011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(667)
);
fnc_OWN668 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010011100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(668)
);
fnc_OWN669 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010011101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(669)
);
fnc_OWN670 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010011110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(670)
);
fnc_OWN671 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010011111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(671)
);
fnc_OWN672 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010100000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(672)
);
fnc_OWN673 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010100001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(673)
);
fnc_OWN674 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010100010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(674)
);
fnc_OWN675 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010100011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(675)
);
fnc_OWN676 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010100100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(676)
);
fnc_OWN677 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010100101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(677)
);
fnc_OWN678 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010100110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(678)
);
fnc_OWN679 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010100111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(679)
);
fnc_OWN680 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010101000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(680)
);
fnc_OWN681 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010101001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(681)
);
fnc_OWN682 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010101010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(682)
);
fnc_OWN683 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010101011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(683)
);
fnc_OWN684 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010101100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(684)
);
fnc_OWN685 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010101101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(685)
);
fnc_OWN686 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010101110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(686)
);
fnc_OWN687 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010101111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(687)
);
fnc_OWN688 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010110000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(688)
);
fnc_OWN689 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010110001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(689)
);
fnc_OWN690 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010110010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(690)
);
fnc_OWN691 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010110011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(691)
);
fnc_OWN692 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010110100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(692)
);
fnc_OWN693 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010110101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(693)
);
fnc_OWN694 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010110110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(694)
);
fnc_OWN695 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010110111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(695)
);
fnc_OWN696 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010111000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(696)
);
fnc_OWN697 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010111001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(697)
);
fnc_OWN698 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010111010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(698)
);
fnc_OWN699 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010111011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(699)
);
fnc_OWN700 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010111100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(700)
);
fnc_OWN701 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010111101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(701)
);
fnc_OWN702 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010111110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(702)
);
fnc_OWN703 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001010111111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(703)
);
fnc_OWN704 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011000000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(704)
);
fnc_OWN705 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011000001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(705)
);
fnc_OWN706 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011000010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(706)
);
fnc_OWN707 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011000011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(707)
);
fnc_OWN708 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011000100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(708)
);
fnc_OWN709 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011000101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(709)
);
fnc_OWN710 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011000110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(710)
);
fnc_OWN711 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011000111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(711)
);
fnc_OWN712 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011001000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(712)
);
fnc_OWN713 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011001001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(713)
);
fnc_OWN714 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011001010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(714)
);
fnc_OWN715 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011001011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(715)
);
fnc_OWN716 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011001100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(716)
);
fnc_OWN717 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011001101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(717)
);
fnc_OWN718 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011001110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(718)
);
fnc_OWN719 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011001111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(719)
);
fnc_OWN720 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011010000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(720)
);
fnc_OWN721 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011010001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(721)
);
fnc_OWN722 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011010010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(722)
);
fnc_OWN723 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011010011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(723)
);
fnc_OWN724 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011010100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(724)
);
fnc_OWN725 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011010101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(725)
);
fnc_OWN726 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011010110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(726)
);
fnc_OWN727 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011010111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(727)
);
fnc_OWN728 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011011000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(728)
);
fnc_OWN729 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011011001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(729)
);
fnc_OWN730 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011011010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(730)
);
fnc_OWN731 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011011011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(731)
);
fnc_OWN732 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011011100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(732)
);
fnc_OWN733 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011011101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(733)
);
fnc_OWN734 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011011110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(734)
);
fnc_OWN735 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011011111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(735)
);
fnc_OWN736 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011100000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(736)
);
fnc_OWN737 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011100001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(737)
);
fnc_OWN738 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011100010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(738)
);
fnc_OWN739 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011100011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(739)
);
fnc_OWN740 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011100100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(740)
);
fnc_OWN741 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011100101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(741)
);
fnc_OWN742 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011100110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(742)
);
fnc_OWN743 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011100111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(743)
);
fnc_OWN744 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011101000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(744)
);
fnc_OWN745 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011101001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(745)
);
fnc_OWN746 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011101010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(746)
);
fnc_OWN747 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011101011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(747)
);
fnc_OWN748 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011101100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(748)
);
fnc_OWN749 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011101101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(749)
);
fnc_OWN750 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011101110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(750)
);
fnc_OWN751 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011101111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(751)
);
fnc_OWN752 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011110000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(752)
);
fnc_OWN753 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011110001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(753)
);
fnc_OWN754 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011110010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(754)
);
fnc_OWN755 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011110011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(755)
);
fnc_OWN756 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011110100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(756)
);
fnc_OWN757 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011110101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(757)
);
fnc_OWN758 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011110110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(758)
);
fnc_OWN759 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011110111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(759)
);
fnc_OWN760 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011111000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(760)
);
fnc_OWN761 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011111001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(761)
);
fnc_OWN762 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011111010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(762)
);
fnc_OWN763 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011111011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(763)
);
fnc_OWN764 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011111100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(764)
);
fnc_OWN765 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011111101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(765)
);
fnc_OWN766 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011111110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(766)
);
fnc_OWN767 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001011111111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(767)
);
fnc_OWN768 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100000000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(768)
);
fnc_OWN769 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100000001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(769)
);
fnc_OWN770 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100000010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(770)
);
fnc_OWN771 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100000011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(771)
);
fnc_OWN772 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100000100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(772)
);
fnc_OWN773 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100000101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(773)
);
fnc_OWN774 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100000110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(774)
);
fnc_OWN775 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100000111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(775)
);
fnc_OWN776 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100001000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(776)
);
fnc_OWN777 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100001001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(777)
);
fnc_OWN778 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100001010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(778)
);
fnc_OWN779 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100001011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(779)
);
fnc_OWN780 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100001100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(780)
);
fnc_OWN781 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100001101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(781)
);
fnc_OWN782 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100001110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(782)
);
fnc_OWN783 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100001111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(783)
);
fnc_OWN784 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100010000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(784)
);
fnc_OWN785 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100010001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(785)
);
fnc_OWN786 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100010010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(786)
);
fnc_OWN787 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100010011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(787)
);
fnc_OWN788 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100010100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(788)
);
fnc_OWN789 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100010101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(789)
);
fnc_OWN790 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100010110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(790)
);
fnc_OWN791 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100010111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(791)
);
fnc_OWN792 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100011000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(792)
);
fnc_OWN793 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100011001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(793)
);
fnc_OWN794 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100011010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(794)
);
fnc_OWN795 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100011011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(795)
);
fnc_OWN796 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100011100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(796)
);
fnc_OWN797 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100011101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(797)
);
fnc_OWN798 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100011110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(798)
);
fnc_OWN799 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100011111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(799)
);
fnc_OWN800 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100100000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(800)
);
fnc_OWN801 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100100001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(801)
);
fnc_OWN802 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100100010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(802)
);
fnc_OWN803 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100100011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(803)
);
fnc_OWN804 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100100100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(804)
);
fnc_OWN805 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100100101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(805)
);
fnc_OWN806 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100100110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(806)
);
fnc_OWN807 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100100111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(807)
);
fnc_OWN808 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100101000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(808)
);
fnc_OWN809 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100101001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(809)
);
fnc_OWN810 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100101010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(810)
);
fnc_OWN811 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100101011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(811)
);
fnc_OWN812 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100101100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(812)
);
fnc_OWN813 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100101101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(813)
);
fnc_OWN814 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100101110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(814)
);
fnc_OWN815 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100101111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(815)
);
fnc_OWN816 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100110000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(816)
);
fnc_OWN817 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100110001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(817)
);
fnc_OWN818 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100110010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(818)
);
fnc_OWN819 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100110011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(819)
);
fnc_OWN820 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100110100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(820)
);
fnc_OWN821 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100110101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(821)
);
fnc_OWN822 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100110110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(822)
);
fnc_OWN823 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100110111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(823)
);
fnc_OWN824 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100111000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(824)
);
fnc_OWN825 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100111001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(825)
);
fnc_OWN826 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100111010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(826)
);
fnc_OWN827 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100111011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(827)
);
fnc_OWN828 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100111100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(828)
);
fnc_OWN829 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100111101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(829)
);
fnc_OWN830 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100111110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(830)
);
fnc_OWN831 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001100111111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(831)
);
fnc_OWN832 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101000000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(832)
);
fnc_OWN833 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101000001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(833)
);
fnc_OWN834 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101000010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(834)
);
fnc_OWN835 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101000011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(835)
);
fnc_OWN836 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101000100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(836)
);
fnc_OWN837 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101000101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(837)
);
fnc_OWN838 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101000110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(838)
);
fnc_OWN839 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101000111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(839)
);
fnc_OWN840 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101001000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(840)
);
fnc_OWN841 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101001001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(841)
);
fnc_OWN842 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101001010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(842)
);
fnc_OWN843 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101001011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(843)
);
fnc_OWN844 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101001100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(844)
);
fnc_OWN845 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101001101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(845)
);
fnc_OWN846 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101001110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(846)
);
fnc_OWN847 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101001111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(847)
);
fnc_OWN848 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101010000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(848)
);
fnc_OWN849 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101010001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(849)
);
fnc_OWN850 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101010010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(850)
);
fnc_OWN851 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101010011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(851)
);
fnc_OWN852 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101010100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(852)
);
fnc_OWN853 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101010101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(853)
);
fnc_OWN854 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101010110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(854)
);
fnc_OWN855 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101010111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(855)
);
fnc_OWN856 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101011000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(856)
);
fnc_OWN857 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101011001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(857)
);
fnc_OWN858 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101011010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(858)
);
fnc_OWN859 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101011011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(859)
);
fnc_OWN860 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101011100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(860)
);
fnc_OWN861 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101011101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(861)
);
fnc_OWN862 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101011110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(862)
);
fnc_OWN863 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101011111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(863)
);
fnc_OWN864 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101100000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(864)
);
fnc_OWN865 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101100001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(865)
);
fnc_OWN866 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101100010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(866)
);
fnc_OWN867 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101100011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(867)
);
fnc_OWN868 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101100100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(868)
);
fnc_OWN869 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101100101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(869)
);
fnc_OWN870 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101100110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(870)
);
fnc_OWN871 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101100111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(871)
);
fnc_OWN872 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101101000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(872)
);
fnc_OWN873 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101101001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(873)
);
fnc_OWN874 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101101010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(874)
);
fnc_OWN875 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101101011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(875)
);
fnc_OWN876 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101101100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(876)
);
fnc_OWN877 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101101101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(877)
);
fnc_OWN878 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101101110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(878)
);
fnc_OWN879 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101101111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(879)
);
fnc_OWN880 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101110000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(880)
);
fnc_OWN881 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101110001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(881)
);
fnc_OWN882 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101110010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(882)
);
fnc_OWN883 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101110011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(883)
);
fnc_OWN884 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101110100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(884)
);
fnc_OWN885 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101110101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(885)
);
fnc_OWN886 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101110110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(886)
);
fnc_OWN887 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101110111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(887)
);
fnc_OWN888 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101111000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(888)
);
fnc_OWN889 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101111001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(889)
);
fnc_OWN890 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101111010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(890)
);
fnc_OWN891 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101111011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(891)
);
fnc_OWN892 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101111100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(892)
);
fnc_OWN893 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101111101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(893)
);
fnc_OWN894 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101111110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(894)
);
fnc_OWN895 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001101111111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(895)
);
fnc_OWN896 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110000000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(896)
);
fnc_OWN897 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110000001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(897)
);
fnc_OWN898 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110000010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(898)
);
fnc_OWN899 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110000011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(899)
);
fnc_OWN900 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110000100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(900)
);
fnc_OWN901 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110000101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(901)
);
fnc_OWN902 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110000110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(902)
);
fnc_OWN903 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110000111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(903)
);
fnc_OWN904 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110001000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(904)
);
fnc_OWN905 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110001001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(905)
);
fnc_OWN906 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110001010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(906)
);
fnc_OWN907 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110001011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(907)
);
fnc_OWN908 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110001100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(908)
);
fnc_OWN909 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110001101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(909)
);
fnc_OWN910 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110001110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(910)
);
fnc_OWN911 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110001111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(911)
);
fnc_OWN912 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110010000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(912)
);
fnc_OWN913 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110010001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(913)
);
fnc_OWN914 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110010010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(914)
);
fnc_OWN915 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110010011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(915)
);
fnc_OWN916 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110010100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(916)
);
fnc_OWN917 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110010101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(917)
);
fnc_OWN918 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110010110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(918)
);
fnc_OWN919 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110010111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(919)
);
fnc_OWN920 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110011000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(920)
);
fnc_OWN921 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110011001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(921)
);
fnc_OWN922 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110011010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(922)
);
fnc_OWN923 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110011011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(923)
);
fnc_OWN924 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110011100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(924)
);
fnc_OWN925 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110011101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(925)
);
fnc_OWN926 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110011110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(926)
);
fnc_OWN927 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110011111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(927)
);
fnc_OWN928 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110100000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(928)
);
fnc_OWN929 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110100001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(929)
);
fnc_OWN930 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110100010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(930)
);
fnc_OWN931 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110100011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(931)
);
fnc_OWN932 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110100100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(932)
);
fnc_OWN933 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110100101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(933)
);
fnc_OWN934 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110100110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(934)
);
fnc_OWN935 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110100111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(935)
);
fnc_OWN936 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110101000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(936)
);
fnc_OWN937 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110101001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(937)
);
fnc_OWN938 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110101010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(938)
);
fnc_OWN939 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110101011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(939)
);
fnc_OWN940 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110101100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(940)
);
fnc_OWN941 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110101101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(941)
);
fnc_OWN942 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110101110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(942)
);
fnc_OWN943 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110101111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(943)
);
fnc_OWN944 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110110000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(944)
);
fnc_OWN945 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110110001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(945)
);
fnc_OWN946 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110110010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(946)
);
fnc_OWN947 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110110011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(947)
);
fnc_OWN948 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110110100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(948)
);
fnc_OWN949 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110110101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(949)
);
fnc_OWN950 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110110110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(950)
);
fnc_OWN951 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110110111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(951)
);
fnc_OWN952 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110111000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(952)
);
fnc_OWN953 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110111001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(953)
);
fnc_OWN954 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110111010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(954)
);
fnc_OWN955 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110111011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(955)
);
fnc_OWN956 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110111100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(956)
);
fnc_OWN957 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110111101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(957)
);
fnc_OWN958 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110111110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(958)
);
fnc_OWN959 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001110111111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(959)
);
fnc_OWN960 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111000000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(960)
);
fnc_OWN961 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111000001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(961)
);
fnc_OWN962 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111000010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(962)
);
fnc_OWN963 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111000011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(963)
);
fnc_OWN964 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111000100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(964)
);
fnc_OWN965 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111000101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(965)
);
fnc_OWN966 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111000110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(966)
);
fnc_OWN967 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111000111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(967)
);
fnc_OWN968 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111001000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(968)
);
fnc_OWN969 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111001001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(969)
);
fnc_OWN970 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111001010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(970)
);
fnc_OWN971 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111001011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(971)
);
fnc_OWN972 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111001100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(972)
);
fnc_OWN973 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111001101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(973)
);
fnc_OWN974 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111001110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(974)
);
fnc_OWN975 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111001111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(975)
);
fnc_OWN976 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111010000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(976)
);
fnc_OWN977 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111010001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(977)
);
fnc_OWN978 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111010010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(978)
);
fnc_OWN979 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111010011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(979)
);
fnc_OWN980 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111010100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(980)
);
fnc_OWN981 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111010101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(981)
);
fnc_OWN982 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111010110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(982)
);
fnc_OWN983 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111010111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(983)
);
fnc_OWN984 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111011000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(984)
);
fnc_OWN985 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111011001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(985)
);
fnc_OWN986 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111011010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(986)
);
fnc_OWN987 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111011011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(987)
);
fnc_OWN988 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111011100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(988)
);
fnc_OWN989 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111011101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(989)
);
fnc_OWN990 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111011110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(990)
);
fnc_OWN991 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111011111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(991)
);
fnc_OWN992 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111100000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(992)
);
fnc_OWN993 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111100001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(993)
);
fnc_OWN994 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111100010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(994)
);
fnc_OWN995 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111100011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(995)
);
fnc_OWN996 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111100100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(996)
);
fnc_OWN997 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111100101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(997)
);
fnc_OWN998 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111100110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(998)
);
fnc_OWN999 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111100111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(999)
);
fnc_OWN1000 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111101000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1000)
);
fnc_OWN1001 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111101001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1001)
);
fnc_OWN1002 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111101010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1002)
);
fnc_OWN1003 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111101011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1003)
);
fnc_OWN1004 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111101100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1004)
);
fnc_OWN1005 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111101101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1005)
);
fnc_OWN1006 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111101110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1006)
);
fnc_OWN1007 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111101111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1007)
);
fnc_OWN1008 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111110000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1008)
);
fnc_OWN1009 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111110001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1009)
);
fnc_OWN1010 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111110010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1010)
);
fnc_OWN1011 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111110011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1011)
);
fnc_OWN1012 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111110100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1012)
);
fnc_OWN1013 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111110101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1013)
);
fnc_OWN1014 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111110110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1014)
);
fnc_OWN1015 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111110111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1015)
);
fnc_OWN1016 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111111000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1016)
);
fnc_OWN1017 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111111001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1017)
);
fnc_OWN1018 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111111010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1018)
);
fnc_OWN1019 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111111011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1019)
);
fnc_OWN1020 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111111100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1020)
);
fnc_OWN1021 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111111101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1021)
);
fnc_OWN1022 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111111110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1022)
);
fnc_OWN1023 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000001111111111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1023)
);
fnc_OWN1024 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000000000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1024)
);
fnc_OWN1025 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000000001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1025)
);
fnc_OWN1026 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000000010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1026)
);
fnc_OWN1027 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000000011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1027)
);
fnc_OWN1028 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000000100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1028)
);
fnc_OWN1029 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000000101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1029)
);
fnc_OWN1030 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000000110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1030)
);
fnc_OWN1031 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000000111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1031)
);
fnc_OWN1032 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000001000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1032)
);
fnc_OWN1033 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000001001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1033)
);
fnc_OWN1034 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000001010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1034)
);
fnc_OWN1035 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000001011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1035)
);
fnc_OWN1036 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000001100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1036)
);
fnc_OWN1037 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000001101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1037)
);
fnc_OWN1038 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000001110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1038)
);
fnc_OWN1039 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000001111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1039)
);
fnc_OWN1040 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000010000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1040)
);
fnc_OWN1041 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000010001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1041)
);
fnc_OWN1042 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000010010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1042)
);
fnc_OWN1043 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000010011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1043)
);
fnc_OWN1044 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000010100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1044)
);
fnc_OWN1045 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000010101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1045)
);
fnc_OWN1046 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000010110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1046)
);
fnc_OWN1047 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000010111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1047)
);
fnc_OWN1048 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000011000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1048)
);
fnc_OWN1049 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000011001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1049)
);
fnc_OWN1050 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000011010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1050)
);
fnc_OWN1051 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000011011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1051)
);
fnc_OWN1052 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000011100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1052)
);
fnc_OWN1053 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000011101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1053)
);
fnc_OWN1054 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000011110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1054)
);
fnc_OWN1055 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000011111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1055)
);
fnc_OWN1056 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000100000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1056)
);
fnc_OWN1057 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000100001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1057)
);
fnc_OWN1058 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000100010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1058)
);
fnc_OWN1059 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000100011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1059)
);
fnc_OWN1060 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000100100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1060)
);
fnc_OWN1061 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000100101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1061)
);
fnc_OWN1062 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000100110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1062)
);
fnc_OWN1063 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000100111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1063)
);
fnc_OWN1064 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000101000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1064)
);
fnc_OWN1065 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000101001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1065)
);
fnc_OWN1066 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000101010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1066)
);
fnc_OWN1067 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000101011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1067)
);
fnc_OWN1068 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000101100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1068)
);
fnc_OWN1069 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000101101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1069)
);
fnc_OWN1070 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000101110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1070)
);
fnc_OWN1071 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000101111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1071)
);
fnc_OWN1072 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000110000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1072)
);
fnc_OWN1073 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000110001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1073)
);
fnc_OWN1074 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000110010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1074)
);
fnc_OWN1075 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000110011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1075)
);
fnc_OWN1076 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000110100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1076)
);
fnc_OWN1077 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000110101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1077)
);
fnc_OWN1078 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000110110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1078)
);
fnc_OWN1079 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000110111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1079)
);
fnc_OWN1080 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000111000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1080)
);
fnc_OWN1081 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000111001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1081)
);
fnc_OWN1082 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000111010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1082)
);
fnc_OWN1083 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000111011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1083)
);
fnc_OWN1084 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000111100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1084)
);
fnc_OWN1085 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000111101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1085)
);
fnc_OWN1086 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000111110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1086)
);
fnc_OWN1087 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010000111111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1087)
);
fnc_OWN1088 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001000000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1088)
);
fnc_OWN1089 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001000001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1089)
);
fnc_OWN1090 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001000010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1090)
);
fnc_OWN1091 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001000011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1091)
);
fnc_OWN1092 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001000100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1092)
);
fnc_OWN1093 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001000101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1093)
);
fnc_OWN1094 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001000110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1094)
);
fnc_OWN1095 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001000111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1095)
);
fnc_OWN1096 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001001000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1096)
);
fnc_OWN1097 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001001001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1097)
);
fnc_OWN1098 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001001010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1098)
);
fnc_OWN1099 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001001011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1099)
);
fnc_OWN1100 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001001100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1100)
);
fnc_OWN1101 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001001101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1101)
);
fnc_OWN1102 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001001110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1102)
);
fnc_OWN1103 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001001111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1103)
);
fnc_OWN1104 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001010000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1104)
);
fnc_OWN1105 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001010001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1105)
);
fnc_OWN1106 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001010010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1106)
);
fnc_OWN1107 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001010011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1107)
);
fnc_OWN1108 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001010100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1108)
);
fnc_OWN1109 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001010101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1109)
);
fnc_OWN1110 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001010110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1110)
);
fnc_OWN1111 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001010111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1111)
);
fnc_OWN1112 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001011000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1112)
);
fnc_OWN1113 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001011001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1113)
);
fnc_OWN1114 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001011010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1114)
);
fnc_OWN1115 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001011011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1115)
);
fnc_OWN1116 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001011100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1116)
);
fnc_OWN1117 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001011101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1117)
);
fnc_OWN1118 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001011110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1118)
);
fnc_OWN1119 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001011111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1119)
);
fnc_OWN1120 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001100000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1120)
);
fnc_OWN1121 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001100001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1121)
);
fnc_OWN1122 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001100010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1122)
);
fnc_OWN1123 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001100011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1123)
);
fnc_OWN1124 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001100100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1124)
);
fnc_OWN1125 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001100101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1125)
);
fnc_OWN1126 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001100110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1126)
);
fnc_OWN1127 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001100111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1127)
);
fnc_OWN1128 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001101000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1128)
);
fnc_OWN1129 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001101001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1129)
);
fnc_OWN1130 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001101010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1130)
);
fnc_OWN1131 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001101011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1131)
);
fnc_OWN1132 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001101100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1132)
);
fnc_OWN1133 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001101101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1133)
);
fnc_OWN1134 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001101110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1134)
);
fnc_OWN1135 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001101111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1135)
);
fnc_OWN1136 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001110000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1136)
);
fnc_OWN1137 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001110001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1137)
);
fnc_OWN1138 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001110010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1138)
);
fnc_OWN1139 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001110011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1139)
);
fnc_OWN1140 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001110100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1140)
);
fnc_OWN1141 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001110101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1141)
);
fnc_OWN1142 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001110110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1142)
);
fnc_OWN1143 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001110111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1143)
);
fnc_OWN1144 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001111000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1144)
);
fnc_OWN1145 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001111001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1145)
);
fnc_OWN1146 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001111010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1146)
);
fnc_OWN1147 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001111011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1147)
);
fnc_OWN1148 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001111100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1148)
);
fnc_OWN1149 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001111101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1149)
);
fnc_OWN1150 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001111110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1150)
);
fnc_OWN1151 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010001111111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1151)
);
fnc_OWN1152 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010000000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1152)
);
fnc_OWN1153 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010000001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1153)
);
fnc_OWN1154 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010000010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1154)
);
fnc_OWN1155 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010000011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1155)
);
fnc_OWN1156 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010000100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1156)
);
fnc_OWN1157 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010000101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1157)
);
fnc_OWN1158 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010000110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1158)
);
fnc_OWN1159 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010000111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1159)
);
fnc_OWN1160 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010001000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1160)
);
fnc_OWN1161 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010001001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1161)
);
fnc_OWN1162 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010001010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1162)
);
fnc_OWN1163 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010001011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1163)
);
fnc_OWN1164 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010001100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1164)
);
fnc_OWN1165 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010001101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1165)
);
fnc_OWN1166 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010001110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1166)
);
fnc_OWN1167 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010001111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1167)
);
fnc_OWN1168 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010010000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1168)
);
fnc_OWN1169 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010010001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1169)
);
fnc_OWN1170 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010010010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1170)
);
fnc_OWN1171 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010010011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1171)
);
fnc_OWN1172 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010010100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1172)
);
fnc_OWN1173 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010010101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1173)
);
fnc_OWN1174 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010010110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1174)
);
fnc_OWN1175 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010010111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1175)
);
fnc_OWN1176 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010011000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1176)
);
fnc_OWN1177 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010011001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1177)
);
fnc_OWN1178 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010011010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1178)
);
fnc_OWN1179 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010011011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1179)
);
fnc_OWN1180 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010011100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1180)
);
fnc_OWN1181 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010011101",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1181)
);
fnc_OWN1182 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010011110",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1182)
);
fnc_OWN1183 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010011111",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1183)
);
fnc_OWN1184 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010100000",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1184)
);
fnc_OWN1185 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010100001",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1185)
);
fnc_OWN1186 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010100010",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1186)
);
fnc_OWN1187 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010100011",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1187)
);
fnc_OWN1188 : matcher generic map (
	G_STRUCTURE         => C_STRCT_SIMPLE,
	G_VALUE_A           => "0000010010100100",
	G_FUNCTION_A        => C_FNCTR_SIMP_SEQ
) port map (
	query_opA_i         => query_i(C_QUERY_OWN),
	match_result_o      => sig_fnc_OWN(1188)
);
bram_APP : xilinx_single_port_ram_no_change generic map (
	RAM_WIDTH => C_BRAM_APP_WIDTH,
	RAM_DEPTH => C_BRAM_APP_DEPTH,
	RAM_PERFORMANCE => "LOW_LATENCY", --"HIGH_PERFORMANCE",
	INIT_FILE => "bram_APP.mem"
) port map (
	clka   => clk_i,
	addra  => query_i(C_QUERY_APP)((clogb2(C_BRAM_APP_DEPTH)-1) downto 0),
	dina   => mem_i(C_BRAM_APP_WIDTH-1 downto 0),
	wea    => meme_i(C_BRAM_APP),
	ena    => '1',
	rsta   => '0',
	regcea => '1',
	douta  => sig_ram_APP
);
fnc_DATE0 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "0001110011101010",
	G_VALUE_B           => "1111000010001111",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(0)
);
fnc_DATE1 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "1011001111100100",
	G_VALUE_B           => "1100001011111011",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(1)
);
fnc_DATE2 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "0010101011011101",
	G_VALUE_B           => "0100100101011101",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(2)
);
fnc_DATE3 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "0000000110101000",
	G_VALUE_B           => "1011010110111111",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(3)
);
fnc_DATE4 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "0001010101000100",
	G_VALUE_B           => "1110011000010100",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(4)
);
fnc_DATE5 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "0011010011110111",
	G_VALUE_B           => "1010110010010011",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(5)
);
fnc_DATE6 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "0000000110011111",
	G_VALUE_B           => "0000010010100110",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(6)
);
fnc_DATE7 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "1101111011010010",
	G_VALUE_B           => "1110111010011001",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(7)
);
fnc_DATE8 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "0001001100000110",
	G_VALUE_B           => "1011111101101000",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(8)
);
fnc_DATE9 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "1110001011011000",
	G_VALUE_B           => "1110011011110100",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(9)
);
fnc_DATE10 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "1011001000110101",
	G_VALUE_B           => "1100110100011000",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(10)
);
fnc_DATE11 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "0010100110011111",
	G_VALUE_B           => "1110100100110000",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(11)
);
fnc_DATE12 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "0010011101001001",
	G_VALUE_B           => "1000100001001111",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(12)
);
fnc_DATE13 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "0011001110101001",
	G_VALUE_B           => "1011001111111010",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(13)
);
fnc_DATE14 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "1010101010111100",
	G_VALUE_B           => "1011110000110100",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(14)
);
fnc_DATE15 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "1000011010110011",
	G_VALUE_B           => "1010000011010100",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(15)
);
fnc_DATE16 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "0001010111001010",
	G_VALUE_B           => "1110000100110110",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(16)
);
fnc_DATE17 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "1000011111101011",
	G_VALUE_B           => "1101100101100011",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(17)
);
fnc_DATE18 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "0001000100001000",
	G_VALUE_B           => "1100101000111111",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(18)
);
fnc_DATE19 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "0000100100000111",
	G_VALUE_B           => "1000011000111001",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(19)
);
fnc_DATE20 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "0101000111110010",
	G_VALUE_B           => "1111001010011110",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(20)
);
fnc_DATE21 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "1001110110011000",
	G_VALUE_B           => "1010111000111111",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(21)
);
fnc_DATE22 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "1001110100000100",
	G_VALUE_B           => "1111100010100100",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(22)
);
fnc_DATE23 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "1000110110000001",
	G_VALUE_B           => "1110000110001000",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(23)
);
fnc_DATE24 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "0100010101110000",
	G_VALUE_B           => "1111011000000100",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(24)
);
fnc_DATE25 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "0100011100011001",
	G_VALUE_B           => "0100110000001010",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(25)
);
fnc_DATE26 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "0010110101100110",
	G_VALUE_B           => "1010001000110000",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(26)
);
fnc_DATE27 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "0010110100001001",
	G_VALUE_B           => "1111100011101111",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(27)
);
fnc_DATE28 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "0010010000011000",
	G_VALUE_B           => "1011000111100100",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(28)
);
fnc_DATE29 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "0110001000001111",
	G_VALUE_B           => "1000010010111001",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(29)
);
fnc_DATE30 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "0000100001001100",
	G_VALUE_B           => "1001000111110101",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(30)
);
fnc_DATE31 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "0001010100000011",
	G_VALUE_B           => "0110000110100000",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(31)
);
fnc_DATE32 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "1010010001111001",
	G_VALUE_B           => "1100110101011000",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(32)
);
fnc_DATE33 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "0001011011110101",
	G_VALUE_B           => "0001110000111100",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(33)
);
fnc_DATE34 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "0110111001110101",
	G_VALUE_B           => "1100001101110010",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(34)
);
fnc_DATE35 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "1001011000010011",
	G_VALUE_B           => "1010110000000111",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(35)
);
fnc_DATE36 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "1001111101001001",
	G_VALUE_B           => "1110000110100110",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(36)
);
fnc_DATE37 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "1000101011101110",
	G_VALUE_B           => "1100101110011011",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(37)
);
fnc_DATE38 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "0101001000000010",
	G_VALUE_B           => "0110011110101001",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(38)
);
fnc_DATE39 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "0110000001000011",
	G_VALUE_B           => "1111010110100110",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(39)
);
fnc_DATE40 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "0111110011011010",
	G_VALUE_B           => "1001011010111010",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(40)
);
fnc_DATE41 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "1110011111010110",
	G_VALUE_B           => "1110100101100100",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(41)
);
fnc_DATE42 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "0011110101110011",
	G_VALUE_B           => "0110110110101001",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(42)
);
fnc_DATE43 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "0110000110011110",
	G_VALUE_B           => "0110111110001000",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(43)
);
fnc_DATE44 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "1110100000101001",
	G_VALUE_B           => "1111001001100001",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(44)
);
fnc_DATE45 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "0010110100011010",
	G_VALUE_B           => "1010110010100000",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(45)
);
fnc_DATE46 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "0011101110001011",
	G_VALUE_B           => "0100011001100010",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(46)
);
fnc_DATE47 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "0101101000100100",
	G_VALUE_B           => "1010010101010101",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(47)
);
fnc_DATE48 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "0001110011010010",
	G_VALUE_B           => "0111000010001010",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(48)
);
fnc_DATE49 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "0000000010110110",
	G_VALUE_B           => "1101110110001001",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(49)
);
fnc_DATE50 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "0000100110100111",
	G_VALUE_B           => "1111011111011010",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(50)
);
fnc_DATE51 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "0010111101011100",
	G_VALUE_B           => "0100110001010110",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(51)
);
fnc_DATE52 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "1010010110100001",
	G_VALUE_B           => "1100101111010001",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(52)
);
fnc_DATE53 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "1010101011101001",
	G_VALUE_B           => "1100011110010111",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(53)
);
fnc_DATE54 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "1001010011110011",
	G_VALUE_B           => "1110011011000111",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(54)
);
fnc_DATE55 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "1000000000000111",
	G_VALUE_B           => "1110111101010000",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(55)
);
fnc_DATE56 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "0010110010001011",
	G_VALUE_B           => "1001001110011111",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(56)
);
fnc_DATE57 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "0100000111010010",
	G_VALUE_B           => "1100100100100110",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(57)
);
fnc_DATE58 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "0010101111000001",
	G_VALUE_B           => "1100010011101110",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(58)
);
fnc_DATE59 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "0101000101111100",
	G_VALUE_B           => "1011100100101010",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(59)
);
fnc_DATE60 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "0011111111010101",
	G_VALUE_B           => "1100001000001100",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(60)
);
fnc_DATE61 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "0001010011100100",
	G_VALUE_B           => "0010000010001000",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(61)
);
fnc_DATE62 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "0000000001110010",
	G_VALUE_B           => "0100000101000001",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(62)
);
fnc_DATE63 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "0100101011110100",
	G_VALUE_B           => "0111011100111110",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(63)
);
fnc_DATE64 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "0110001100100101",
	G_VALUE_B           => "1111101010110111",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(64)
);
fnc_DATE65 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "1011010110101110",
	G_VALUE_B           => "1100011010000101",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(65)
);
fnc_DATE66 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "0110000010001011",
	G_VALUE_B           => "1010001111111101",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(66)
);
fnc_DATE67 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "1000100001111101",
	G_VALUE_B           => "1010010101110111",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(67)
);
fnc_DATE68 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "0001111001110010",
	G_VALUE_B           => "0101111100110001",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(68)
);
fnc_DATE69 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "0001011101001011",
	G_VALUE_B           => "0001100001111001",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(69)
);
fnc_DATE70 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "0110011001010100",
	G_VALUE_B           => "1100101011011110",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(70)
);
fnc_DATE71 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "1000001010000101",
	G_VALUE_B           => "1110000100100101",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(71)
);
fnc_DATE72 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "0011100100111000",
	G_VALUE_B           => "1100100011010010",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(72)
);
fnc_DATE73 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "0101010010110110",
	G_VALUE_B           => "1111101110111100",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(73)
);
fnc_DATE74 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "0011100101011100",
	G_VALUE_B           => "1011100001011001",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(74)
);
fnc_DATE75 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "0001111011010110",
	G_VALUE_B           => "1111111101111010",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(75)
);
fnc_DATE76 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "1000100010110000",
	G_VALUE_B           => "1010001000010100",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(76)
);
fnc_DATE77 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "0111001110011000",
	G_VALUE_B           => "1000111010010110",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(77)
);
fnc_DATE78 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "0001101011000111",
	G_VALUE_B           => "0110000011101010",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(78)
);
fnc_DATE79 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "0101011101111001",
	G_VALUE_B           => "1011011011011101",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(79)
);
fnc_DATE80 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "0010111010110111",
	G_VALUE_B           => "1111010111100101",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(80)
);
fnc_DATE81 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "0001111111011110",
	G_VALUE_B           => "0011001011100101",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(81)
);
fnc_DATE82 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "0100001111111000",
	G_VALUE_B           => "1000010011101111",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(82)
);
fnc_DATE83 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "0001001010001000",
	G_VALUE_B           => "0101111111001100",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(83)
);
fnc_DATE84 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "1101100011111001",
	G_VALUE_B           => "1110001101011111",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(84)
);
fnc_DATE85 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "0000000001011011",
	G_VALUE_B           => "1011011110101111",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(85)
);
fnc_DATE86 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "0010110001110001",
	G_VALUE_B           => "1011110001111110",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(86)
);
fnc_DATE87 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "0000001011000100",
	G_VALUE_B           => "1010000011100111",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(87)
);
fnc_DATE88 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "0101001000111101",
	G_VALUE_B           => "1000000101011100",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(88)
);
fnc_DATE89 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "0101111000110111",
	G_VALUE_B           => "1011001101001101",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(89)
);
fnc_DATE90 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "0010000101000001",
	G_VALUE_B           => "0100100110011010",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(90)
);
fnc_DATE91 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "1100111000100000",
	G_VALUE_B           => "1101011110110101",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(91)
);
fnc_DATE92 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "0110100100101101",
	G_VALUE_B           => "0111010011101011",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(92)
);
fnc_DATE93 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "0110110011110000",
	G_VALUE_B           => "1111110000010101",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(93)
);
fnc_DATE94 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "0111000010001101",
	G_VALUE_B           => "0111111111001111",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(94)
);
fnc_DATE95 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "0001001010000010",
	G_VALUE_B           => "1111001110110100",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(95)
);
fnc_DATE96 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "0100110111001011",
	G_VALUE_B           => "0110010011000011",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(96)
);
fnc_DATE97 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "0110000000011001",
	G_VALUE_B           => "1100110001100000",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(97)
);
fnc_DATE98 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "0111111100111011",
	G_VALUE_B           => "1110011100011111",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(98)
);
fnc_DATE99 : matcher generic map (
	G_STRUCTURE         => C_STRCT_PAIR,
	G_VALUE_A           => "0011100010100110",
	G_VALUE_B           => "0110011101110001",
	G_FUNCTION_A        => C_FNCTR_SIMP_DSE,
	G_FUNCTION_B        => C_FNCTR_SIMP_DIE,
	G_FUNCTION_PAIR     => C_FNCTR_PAIR_PCA
) port map (
	query_opA_i         => query_i(C_QUERY_DATEA),
	query_opB_i         => query_i(C_QUERY_DATEB),
	match_result_o      => sig_fnc_DATE(99)
);
bram_MKTA : xilinx_single_port_ram_no_change generic map (
	RAM_WIDTH => C_BRAM_MKTA_WIDTH,
	RAM_DEPTH => C_BRAM_MKTA_DEPTH,
	RAM_PERFORMANCE => "LOW_LATENCY", --"HIGH_PERFORMANCE",
	INIT_FILE => "bram_MKTA.mem"
) port map (
	clka   => clk_i,
	addra  => query_i(C_QUERY_MKTA)((clogb2(C_BRAM_MKTA_DEPTH)-1) downto 0),
	dina   => mem_i(C_BRAM_MKTA_WIDTH-1 downto 0),
	wea    => meme_i(C_BRAM_MKTA),
	ena    => '1',
	rsta   => '0',
	regcea => '1',
	douta  => sig_ram_MKTA
);
bram_MKTB : xilinx_single_port_ram_no_change generic map (
	RAM_WIDTH => C_BRAM_MKTB_WIDTH,
	RAM_DEPTH => C_BRAM_MKTB_DEPTH,
	RAM_PERFORMANCE => "LOW_LATENCY", --"HIGH_PERFORMANCE",
	INIT_FILE => "bram_MKTB.mem"
) port map (
	clka   => clk_i,
	addra  => query_i(C_QUERY_MKTB)((clogb2(C_BRAM_MKTB_DEPTH)-1) downto 0),
	dina   => mem_i(C_BRAM_MKTB_WIDTH-1 downto 0),
	wea    => meme_i(C_BRAM_MKTB),
	ena    => '1',
	rsta   => '0',
	regcea => '1',
	douta  => sig_ram_MKTB
);
bram_CABIN : xilinx_single_port_ram_no_change generic map (
	RAM_WIDTH => C_BRAM_CABIN_WIDTH,
	RAM_DEPTH => C_BRAM_CABIN_DEPTH,
	RAM_PERFORMANCE => "LOW_LATENCY", --"HIGH_PERFORMANCE",
	INIT_FILE => "bram_CABIN.mem"
) port map (
	clka   => clk_i,
	addra  => query_i(C_QUERY_CABIN)((clogb2(C_BRAM_CABIN_DEPTH)-1) downto 0),
	dina   => mem_i(C_BRAM_CABIN_WIDTH-1 downto 0),
	wea    => meme_i(C_BRAM_CABIN),
	ena    => '1',
	rsta   => '0',
	regcea => '1',
	douta  => sig_ram_CABIN
);
bram_BKG : xilinx_single_port_ram_no_change generic map (
	RAM_WIDTH => C_BRAM_BKG_WIDTH,
	RAM_DEPTH => C_BRAM_BKG_DEPTH,
	RAM_PERFORMANCE => "LOW_LATENCY", --"HIGH_PERFORMANCE",
	INIT_FILE => "bram_BKG.mem"
) port map (
	clka   => clk_i,
	addra  => query_i(C_QUERY_BKG)((clogb2(C_BRAM_BKG_DEPTH)-1) downto 0),
	dina   => mem_i(C_BRAM_BKG_WIDTH-1 downto 0),
	wea    => meme_i(C_BRAM_BKG),
	ena    => '1',
	rsta   => '0',
	regcea => '1',
	douta  => sig_ram_BKG
);
sig_rule(0000000) <= 
		sig_fnc_RTD(1582)
		sig_ram_VERS(4)
		sig_fnc_OWN(709)
		sig_ram_APP(23)
		sig_fnc_DATE(60)
		sig_ram_MKTA(2)
		sig_ram_MKTB(23)
		sig_ram_CABIN(2)
		sig_ram_BKG(3);
sig_rule(0000001) <= 
		sig_fnc_RTD(2080)
		sig_ram_VERS(4)
		sig_fnc_OWN(946)
		sig_ram_APP(10)
		sig_fnc_DATE(9)
		sig_ram_MKTA(15)
		sig_ram_MKTB(22)
		sig_ram_CABIN(3)
		sig_ram_BKG(19);
sig_rule(0000002) <= 
		sig_fnc_RTD(1840)
		sig_ram_VERS(3)
		sig_fnc_OWN(296)
		sig_ram_APP(12)
		sig_fnc_DATE(37)
		sig_ram_MKTA(21)
		sig_ram_MKTB(4)
		sig_ram_CABIN(1)
		sig_ram_BKG(1);
sig_rule(0000003) <= 
		sig_fnc_RTD(1058)
		sig_ram_VERS(4)
		sig_fnc_OWN(798)
		sig_ram_APP(24)
		sig_fnc_DATE(67)
		sig_ram_MKTA(7)
		sig_ram_MKTB(17)
		sig_ram_CABIN(7)
		sig_ram_BKG(12);
sig_rule(0000004) <= 
		sig_fnc_RTD(728)
		sig_ram_VERS(3)
		sig_fnc_OWN(365)
		sig_ram_APP(32)
		sig_fnc_DATE(43)
		sig_ram_MKTA(0);
sig_rule(0000005) <= 
		sig_fnc_RTD(1889)
		sig_ram_VERS(4)
		sig_fnc_OWN(506)
		sig_ram_APP(2)
		sig_fnc_DATE(55)
		sig_ram_MKTA(22)
		sig_ram_MKTB(26)
		sig_ram_CABIN(2)
		sig_ram_BKG(17);
sig_rule(0000006) <= 
		sig_fnc_RTD(2004)
		sig_ram_VERS(0)
		sig_fnc_OWN(1185)
		sig_ram_APP(23)
		sig_fnc_DATE(43)
		sig_ram_MKTA(31)
		sig_ram_MKTB(26)
		sig_ram_CABIN(5)
		sig_ram_BKG(1);
sig_rule(0000007) <= 
		sig_fnc_RTD(1594)
		sig_ram_VERS(1)
		sig_fnc_OWN(153)
		sig_ram_APP(6)
		sig_fnc_DATE(70)
		sig_ram_MKTA(23)
		sig_ram_MKTB(14)
		sig_ram_CABIN(1)
		sig_ram_BKG(1);
sig_rule(0000008) <= 
		sig_fnc_RTD(484)
		sig_ram_VERS(1)
		sig_fnc_OWN(665)
		sig_ram_APP(15)
		sig_fnc_DATE(7)
		sig_ram_MKTA(4)
		sig_ram_MKTB(4)
		sig_ram_CABIN(2)
		sig_ram_BKG(8);
sig_rule(0000009) <= 
		sig_fnc_RTD(1759)
		sig_ram_VERS(0)
		sig_fnc_OWN(542)
		sig_ram_APP(8)
		sig_fnc_DATE(4)
		sig_ram_MKTA(18)
		sig_ram_MKTB(31)
		sig_ram_CABIN(4)
		sig_ram_BKG(16);
sig_rule(0000010) <= 
		sig_fnc_RTD(842)
		sig_ram_VERS(1)
		sig_fnc_OWN(80)
		sig_ram_APP(32)
		sig_fnc_DATE(31)
		sig_ram_MKTA(1)
		sig_ram_MKTB(17)
		sig_ram_CABIN(6)
		sig_ram_BKG(10);
sig_rule(0000011) <= 
		sig_fnc_RTD(375)
		sig_ram_VERS(4)
		sig_fnc_OWN(809)
		sig_ram_APP(20)
		sig_fnc_DATE(88)
		sig_ram_MKTA(28)
		sig_ram_MKTB(14)
		sig_ram_CABIN(0);
sig_rule(0000012) <= 
		sig_fnc_RTD(2701)
		sig_ram_VERS(1)
		sig_fnc_OWN(75)
		sig_ram_APP(22)
		sig_fnc_DATE(29)
		sig_ram_MKTA(11)
		sig_ram_MKTB(26)
		sig_ram_CABIN(0);
sig_rule(0000013) <= 
		sig_fnc_RTD(519)
		sig_ram_VERS(4)
		sig_fnc_OWN(942)
		sig_ram_APP(31)
		sig_fnc_DATE(60)
		sig_ram_MKTA(26)
		sig_ram_MKTB(25)
		sig_ram_CABIN(2)
		sig_ram_BKG(13);
sig_rule(0000014) <= 
		sig_fnc_RTD(2410)
		sig_ram_VERS(0)
		sig_fnc_OWN(484)
		sig_ram_APP(37)
		sig_fnc_DATE(59)
		sig_ram_MKTA(24)
		sig_ram_MKTB(26)
		sig_ram_CABIN(6)
		sig_ram_BKG(1);
sig_rule(0000015) <= 
		sig_fnc_RTD(1036)
		sig_ram_VERS(1)
		sig_fnc_OWN(11)
		sig_ram_APP(25)
		sig_fnc_DATE(68)
		sig_ram_MKTA(4)
		sig_ram_MKTB(13)
		sig_ram_CABIN(1)
		sig_ram_BKG(10);
sig_rule(0000016) <= 
		sig_fnc_RTD(593)
		sig_ram_VERS(3)
		sig_fnc_OWN(248)
		sig_ram_APP(44)
		sig_fnc_DATE(22)
		sig_ram_MKTA(14)
		sig_ram_MKTB(12)
		sig_ram_CABIN(0);
sig_rule(0000017) <= 
		sig_fnc_RTD(261)
		sig_ram_VERS(4)
		sig_fnc_OWN(776)
		sig_ram_APP(32)
		sig_fnc_DATE(61)
		sig_ram_MKTA(6)
		sig_ram_MKTB(23)
		sig_ram_CABIN(0);
sig_rule(0000018) <= 
		sig_fnc_RTD(1362)
		sig_ram_VERS(2)
		sig_fnc_OWN(1175)
		sig_ram_APP(27)
		sig_fnc_DATE(4)
		sig_ram_MKTA(7)
		sig_ram_MKTB(0);
sig_rule(0000019) <= 
		sig_fnc_RTD(2667)
		sig_ram_VERS(2)
		sig_fnc_OWN(254)
		sig_ram_APP(19)
		sig_fnc_DATE(19)
		sig_ram_MKTA(31)
		sig_ram_MKTB(27)
		sig_ram_CABIN(2)
		sig_ram_BKG(9);
sig_rule(0000020) <= 
		sig_fnc_RTD(1689)
		sig_ram_VERS(2)
		sig_fnc_OWN(742)
		sig_ram_APP(30)
		sig_fnc_DATE(20)
		sig_ram_MKTA(0);
sig_rule(0000021) <= 
		sig_fnc_RTD(1015)
		sig_ram_VERS(4)
		sig_fnc_OWN(891)
		sig_ram_APP(24)
		sig_fnc_DATE(27)
		sig_ram_MKTA(27)
		sig_ram_MKTB(2)
		sig_ram_CABIN(0);
sig_rule(0000022) <= 
		sig_fnc_RTD(577)
		sig_ram_VERS(3)
		sig_fnc_OWN(648)
		sig_ram_APP(36)
		sig_fnc_DATE(51)
		sig_ram_MKTA(23)
		sig_ram_MKTB(15)
		sig_ram_CABIN(4)
		sig_ram_BKG(14);
sig_rule(0000023) <= 
		sig_fnc_RTD(2240)
		sig_ram_VERS(0)
		sig_fnc_OWN(609)
		sig_ram_APP(36)
		sig_fnc_DATE(3)
		sig_ram_MKTA(2)
		sig_ram_MKTB(9)
		sig_ram_CABIN(5)
		sig_ram_BKG(4);
sig_rule(0000024) <= 
		sig_fnc_RTD(2388)
		sig_ram_VERS(2)
		sig_fnc_OWN(660)
		sig_ram_APP(8)
		sig_fnc_DATE(51)
		sig_ram_MKTA(26)
		sig_ram_MKTB(22)
		sig_ram_CABIN(3)
		sig_ram_BKG(10);
sig_rule(0000025) <= 
		sig_fnc_RTD(982)
		sig_ram_VERS(1)
		sig_fnc_OWN(672)
		sig_ram_APP(35)
		sig_fnc_DATE(69)
		sig_ram_MKTA(22)
		sig_ram_MKTB(8)
		sig_ram_CABIN(3)
		sig_ram_BKG(17);
sig_rule(0000026) <= 
		sig_fnc_RTD(1834)
		sig_ram_VERS(0)
		sig_fnc_OWN(219)
		sig_ram_APP(43)
		sig_fnc_DATE(63)
		sig_ram_MKTA(10)
		sig_ram_MKTB(2)
		sig_ram_CABIN(1)
		sig_ram_BKG(10);
sig_rule(0000027) <= 
		sig_fnc_RTD(1442)
		sig_ram_VERS(1)
		sig_fnc_OWN(579)
		sig_ram_APP(36)
		sig_fnc_DATE(9)
		sig_ram_MKTA(24)
		sig_ram_MKTB(26)
		sig_ram_CABIN(2)
		sig_ram_BKG(1);
sig_rule(0000028) <= 
		sig_fnc_RTD(1846)
		sig_ram_VERS(1)
		sig_fnc_OWN(870)
		sig_ram_APP(27)
		sig_fnc_DATE(67)
		sig_ram_MKTA(2)
		sig_ram_MKTB(16)
		sig_ram_CABIN(7)
		sig_ram_BKG(12);
sig_rule(0000029) <= 
		sig_fnc_RTD(1745)
		sig_ram_VERS(0)
		sig_fnc_OWN(66)
		sig_ram_APP(25)
		sig_fnc_DATE(2)
		sig_ram_MKTA(13)
		sig_ram_MKTB(21)
		sig_ram_CABIN(7)
		sig_ram_BKG(11);
sig_rule(0000030) <= 
		sig_fnc_RTD(2474)
		sig_ram_VERS(0)
		sig_fnc_OWN(952)
		sig_ram_APP(32)
		sig_fnc_DATE(84)
		sig_ram_MKTA(26)
		sig_ram_MKTB(29)
		sig_ram_CABIN(7)
		sig_ram_BKG(25);
sig_rule(0000031) <= 
		sig_fnc_RTD(1933)
		sig_ram_VERS(0)
		sig_fnc_OWN(27)
		sig_ram_APP(44)
		sig_fnc_DATE(11)
		sig_ram_MKTA(1)
		sig_ram_MKTB(10)
		sig_ram_CABIN(7)
		sig_ram_BKG(1);
sig_rule(0000032) <= 
		sig_fnc_RTD(256)
		sig_ram_VERS(4)
		sig_fnc_OWN(634)
		sig_ram_APP(39)
		sig_fnc_DATE(90)
		sig_ram_MKTA(26)
		sig_ram_MKTB(24)
		sig_ram_CABIN(1)
		sig_ram_BKG(14);
sig_rule(0000033) <= 
		sig_fnc_RTD(595)
		sig_ram_VERS(1)
		sig_fnc_OWN(373)
		sig_ram_APP(0);
sig_rule(0000034) <= 
		sig_fnc_RTD(931)
		sig_ram_VERS(1)
		sig_fnc_OWN(313)
		sig_ram_APP(16)
		sig_fnc_DATE(54)
		sig_ram_MKTA(6)
		sig_ram_MKTB(10)
		sig_ram_CABIN(2)
		sig_ram_BKG(7);
sig_rule(0000035) <= 
		sig_fnc_RTD(826)
		sig_ram_VERS(1)
		sig_fnc_OWN(376)
		sig_ram_APP(33)
		sig_fnc_DATE(42)
		sig_ram_MKTA(27)
		sig_ram_MKTB(0);
sig_rule(0000036) <= 
		sig_fnc_RTD(2452)
		sig_ram_VERS(1)
		sig_fnc_OWN(1106)
		sig_ram_APP(34)
		sig_fnc_DATE(64)
		sig_ram_MKTA(19)
		sig_ram_MKTB(8)
		sig_ram_CABIN(3)
		sig_ram_BKG(10);
sig_rule(0000037) <= 
		sig_fnc_RTD(557)
		sig_ram_VERS(3)
		sig_fnc_OWN(901)
		sig_ram_APP(9)
		sig_fnc_DATE(7)
		sig_ram_MKTA(0);
sig_rule(0000038) <= 
		sig_fnc_RTD(2606)
		sig_ram_VERS(0)
		sig_fnc_OWN(808)
		sig_ram_APP(37)
		sig_fnc_DATE(99)
		sig_ram_MKTA(24)
		sig_ram_MKTB(3)
		sig_ram_CABIN(5)
		sig_ram_BKG(20);
sig_rule(0000039) <= 
		sig_fnc_RTD(672)
		sig_ram_VERS(4)
		sig_fnc_OWN(901)
		sig_ram_APP(36)
		sig_fnc_DATE(97)
		sig_ram_MKTA(23)
		sig_ram_MKTB(16)
		sig_ram_CABIN(0);
sig_rule(0000040) <= 
		sig_fnc_RTD(164)
		sig_ram_VERS(4)
		sig_fnc_OWN(709)
		sig_ram_APP(39)
		sig_fnc_DATE(97)
		sig_ram_MKTA(4)
		sig_ram_MKTB(19)
		sig_ram_CABIN(6)
		sig_ram_BKG(15);
sig_rule(0000041) <= 
		sig_fnc_RTD(2776)
		sig_ram_VERS(2)
		sig_fnc_OWN(375)
		sig_ram_APP(10)
		sig_fnc_DATE(54)
		sig_ram_MKTA(27)
		sig_ram_MKTB(19)
		sig_ram_CABIN(0);
sig_rule(0000042) <= 
		sig_fnc_RTD(1575)
		sig_ram_VERS(3)
		sig_fnc_OWN(100)
		sig_ram_APP(3)
		sig_fnc_DATE(62)
		sig_ram_MKTA(5)
		sig_ram_MKTB(16)
		sig_ram_CABIN(0);
sig_rule(0000043) <= 
		sig_fnc_RTD(1149)
		sig_ram_VERS(3)
		sig_fnc_OWN(1040)
		sig_ram_APP(26)
		sig_fnc_DATE(38)
		sig_ram_MKTA(7)
		sig_ram_MKTB(6)
		sig_ram_CABIN(0);
sig_rule(0000044) <= 
		sig_fnc_RTD(159)
		sig_ram_VERS(2)
		sig_fnc_OWN(714)
		sig_ram_APP(35)
		sig_fnc_DATE(84)
		sig_ram_MKTA(10)
		sig_ram_MKTB(0);
sig_rule(0000045) <= 
		sig_fnc_RTD(2650)
		sig_ram_VERS(2)
		sig_fnc_OWN(468)
		sig_ram_APP(5)
		sig_fnc_DATE(69)
		sig_ram_MKTA(1)
		sig_ram_MKTB(22)
		sig_ram_CABIN(1)
		sig_ram_BKG(18);
sig_rule(0000046) <= 
		sig_fnc_RTD(1032)
		sig_ram_VERS(4)
		sig_fnc_OWN(457)
		sig_ram_APP(41)
		sig_fnc_DATE(47)
		sig_ram_MKTA(30)
		sig_ram_MKTB(25)
		sig_ram_CABIN(4)
		sig_ram_BKG(7);
sig_rule(0000047) <= 
		sig_fnc_RTD(251)
		sig_ram_VERS(0)
		sig_fnc_OWN(75)
		sig_ram_APP(39)
		sig_fnc_DATE(38)
		sig_ram_MKTA(16)
		sig_ram_MKTB(13)
		sig_ram_CABIN(4)
		sig_ram_BKG(24);
sig_rule(0000048) <= 
		sig_fnc_RTD(1410)
		sig_ram_VERS(4)
		sig_fnc_OWN(482)
		sig_ram_APP(41)
		sig_fnc_DATE(15)
		sig_ram_MKTA(4)
		sig_ram_MKTB(20)
		sig_ram_CABIN(1)
		sig_ram_BKG(13);
sig_rule(0000049) <= 
		sig_fnc_RTD(772)
		sig_ram_VERS(3)
		sig_fnc_OWN(478)
		sig_ram_APP(10)
		sig_fnc_DATE(81)
		sig_ram_MKTA(26)
		sig_ram_MKTB(26)
		sig_ram_CABIN(3)
		sig_ram_BKG(17);
sig_rule(0000050) <= 
		sig_fnc_RTD(317)
		sig_ram_VERS(3)
		sig_fnc_OWN(1087)
		sig_ram_APP(27)
		sig_fnc_DATE(8)
		sig_ram_MKTA(25)
		sig_ram_MKTB(14)
		sig_ram_CABIN(1)
		sig_ram_BKG(9);
sig_rule(0000051) <= 
		sig_fnc_RTD(1886)
		sig_ram_VERS(4)
		sig_fnc_OWN(1010)
		sig_ram_APP(19)
		sig_fnc_DATE(27)
		sig_ram_MKTA(6)
		sig_ram_MKTB(24)
		sig_ram_CABIN(5)
		sig_ram_BKG(2);
sig_rule(0000052) <= 
		sig_fnc_RTD(1572)
		sig_ram_VERS(2)
		sig_fnc_OWN(459)
		sig_ram_APP(11)
		sig_fnc_DATE(55)
		sig_ram_MKTA(24)
		sig_ram_MKTB(19)
		sig_ram_CABIN(7)
		sig_ram_BKG(12);
sig_rule(0000053) <= 
		sig_fnc_RTD(1743)
		sig_ram_VERS(4)
		sig_fnc_OWN(1095)
		sig_ram_APP(15)
		sig_fnc_DATE(69)
		sig_ram_MKTA(0);
sig_rule(0000054) <= 
		sig_fnc_RTD(1530)
		sig_ram_VERS(2)
		sig_fnc_OWN(522)
		sig_ram_APP(1)
		sig_fnc_DATE(68)
		sig_ram_MKTA(29)
		sig_ram_MKTB(26)
		sig_ram_CABIN(0);
sig_rule(0000055) <= 
		sig_fnc_RTD(70)
		sig_ram_VERS(0)
		sig_fnc_OWN(232)
		sig_ram_APP(2)
		sig_fnc_DATE(84)
		sig_ram_MKTA(10)
		sig_ram_MKTB(12)
		sig_ram_CABIN(4)
		sig_ram_BKG(5);
sig_rule(0000056) <= 
		sig_fnc_RTD(1689)
		sig_ram_VERS(1)
		sig_fnc_OWN(701)
		sig_ram_APP(3)
		sig_fnc_DATE(81)
		sig_ram_MKTA(4)
		sig_ram_MKTB(13)
		sig_ram_CABIN(2)
		sig_ram_BKG(4);
sig_rule(0000057) <= 
		sig_fnc_RTD(2640)
		sig_ram_VERS(4)
		sig_fnc_OWN(1072)
		sig_ram_APP(27)
		sig_fnc_DATE(0);
sig_rule(0000058) <= 
		sig_fnc_RTD(2122)
		sig_ram_VERS(2)
		sig_fnc_OWN(221)
		sig_ram_APP(29)
		sig_fnc_DATE(11)
		sig_ram_MKTA(28)
		sig_ram_MKTB(20)
		sig_ram_CABIN(0);
sig_rule(0000059) <= 
		sig_fnc_RTD(1775)
		sig_ram_VERS(0)
		sig_fnc_OWN(481)
		sig_ram_APP(7)
		sig_fnc_DATE(92)
		sig_ram_MKTA(18)
		sig_ram_MKTB(3)
		sig_ram_CABIN(7)
		sig_ram_BKG(11);
sig_rule(0000060) <= 
		sig_fnc_RTD(2430)
		sig_ram_VERS(2)
		sig_fnc_OWN(394)
		sig_ram_APP(14)
		sig_fnc_DATE(18)
		sig_ram_MKTA(31)
		sig_ram_MKTB(8)
		sig_ram_CABIN(3)
		sig_ram_BKG(20);
sig_rule(0000061) <= 
		sig_fnc_RTD(2395)
		sig_ram_VERS(3)
		sig_fnc_OWN(294)
		sig_ram_APP(33)
		sig_fnc_DATE(5)
		sig_ram_MKTA(18)
		sig_ram_MKTB(10)
		sig_ram_CABIN(5)
		sig_ram_BKG(12);
sig_rule(0000062) <= 
		sig_fnc_RTD(1057)
		sig_ram_VERS(3)
		sig_fnc_OWN(700)
		sig_ram_APP(31)
		sig_fnc_DATE(29)
		sig_ram_MKTA(18)
		sig_ram_MKTB(21)
		sig_ram_CABIN(7)
		sig_ram_BKG(18);
sig_rule(0000063) <= 
		sig_fnc_RTD(1958)
		sig_ram_VERS(2)
		sig_fnc_OWN(514)
		sig_ram_APP(27)
		sig_fnc_DATE(27)
		sig_ram_MKTA(0);
sig_rule(0000064) <= 
		sig_fnc_RTD(1643)
		sig_ram_VERS(3)
		sig_fnc_OWN(918)
		sig_ram_APP(23)
		sig_fnc_DATE(14)
		sig_ram_MKTA(28)
		sig_ram_MKTB(20)
		sig_ram_CABIN(2)
		sig_ram_BKG(2);
sig_rule(0000065) <= 
		sig_fnc_RTD(902)
		sig_ram_VERS(0)
		sig_fnc_OWN(233)
		sig_ram_APP(4)
		sig_fnc_DATE(91)
		sig_ram_MKTA(5)
		sig_ram_MKTB(31)
		sig_ram_CABIN(3)
		sig_ram_BKG(9);
sig_rule(0000066) <= 
		sig_fnc_RTD(937)
		sig_ram_VERS(4)
		sig_fnc_OWN(1084)
		sig_ram_APP(42)
		sig_fnc_DATE(58)
		sig_ram_MKTA(30)
		sig_ram_MKTB(6)
		sig_ram_CABIN(3)
		sig_ram_BKG(24);
sig_rule(0000067) <= 
		sig_fnc_RTD(1972)
		sig_ram_VERS(3)
		sig_fnc_OWN(435)
		sig_ram_APP(5)
		sig_fnc_DATE(59)
		sig_ram_MKTA(18)
		sig_ram_MKTB(21)
		sig_ram_CABIN(6)
		sig_ram_BKG(10);
sig_rule(0000068) <= 
		sig_fnc_RTD(764)
		sig_ram_VERS(4)
		sig_fnc_OWN(846)
		sig_ram_APP(29)
		sig_fnc_DATE(87)
		sig_ram_MKTA(1)
		sig_ram_MKTB(3)
		sig_ram_CABIN(3)
		sig_ram_BKG(20);
sig_rule(0000069) <= 
		sig_fnc_RTD(1665)
		sig_ram_VERS(0)
		sig_fnc_OWN(452)
		sig_ram_APP(9)
		sig_fnc_DATE(77)
		sig_ram_MKTA(21)
		sig_ram_MKTB(17)
		sig_ram_CABIN(7)
		sig_ram_BKG(20);
sig_rule(0000070) <= 
		sig_fnc_RTD(1029)
		sig_ram_VERS(2)
		sig_fnc_OWN(624)
		sig_ram_APP(38)
		sig_fnc_DATE(76)
		sig_ram_MKTA(21)
		sig_ram_MKTB(13)
		sig_ram_CABIN(6)
		sig_ram_BKG(23);
sig_rule(0000071) <= 
		sig_fnc_RTD(1790)
		sig_ram_VERS(2)
		sig_fnc_OWN(212)
		sig_ram_APP(15)
		sig_fnc_DATE(95)
		sig_ram_MKTA(17)
		sig_ram_MKTB(8)
		sig_ram_CABIN(2)
		sig_ram_BKG(8);
sig_rule(0000072) <= 
		sig_fnc_RTD(114)
		sig_ram_VERS(0)
		sig_fnc_OWN(1084)
		sig_ram_APP(14)
		sig_fnc_DATE(28)
		sig_ram_MKTA(9)
		sig_ram_MKTB(8)
		sig_ram_CABIN(1)
		sig_ram_BKG(18);
sig_rule(0000073) <= 
		sig_fnc_RTD(2534)
		sig_ram_VERS(3)
		sig_fnc_OWN(491)
		sig_ram_APP(2)
		sig_fnc_DATE(26)
		sig_ram_MKTA(7)
		sig_ram_MKTB(20)
		sig_ram_CABIN(5)
		sig_ram_BKG(1);
sig_rule(0000074) <= 
		sig_fnc_RTD(1120)
		sig_ram_VERS(1)
		sig_fnc_OWN(229)
		sig_ram_APP(29)
		sig_fnc_DATE(67)
		sig_ram_MKTA(16)
		sig_ram_MKTB(16)
		sig_ram_CABIN(0);
sig_rule(0000075) <= 
		sig_fnc_RTD(1832)
		sig_ram_VERS(1)
		sig_fnc_OWN(650)
		sig_ram_APP(44)
		sig_fnc_DATE(83)
		sig_ram_MKTA(5)
		sig_ram_MKTB(3)
		sig_ram_CABIN(7)
		sig_ram_BKG(5);
sig_rule(0000076) <= 
		sig_fnc_RTD(492)
		sig_ram_VERS(2)
		sig_fnc_OWN(358)
		sig_ram_APP(35)
		sig_fnc_DATE(77)
		sig_ram_MKTA(1)
		sig_ram_MKTB(11)
		sig_ram_CABIN(4)
		sig_ram_BKG(16);
sig_rule(0000077) <= 
		sig_fnc_RTD(1446)
		sig_ram_VERS(4)
		sig_fnc_OWN(43)
		sig_ram_APP(23)
		sig_fnc_DATE(72)
		sig_ram_MKTA(27)
		sig_ram_MKTB(8)
		sig_ram_CABIN(6)
		sig_ram_BKG(7);
sig_rule(0000078) <= 
		sig_fnc_RTD(1566)
		sig_ram_VERS(4)
		sig_fnc_OWN(786)
		sig_ram_APP(10)
		sig_fnc_DATE(12)
		sig_ram_MKTA(8)
		sig_ram_MKTB(14)
		sig_ram_CABIN(3)
		sig_ram_BKG(5);
sig_rule(0000079) <= 
		sig_fnc_RTD(2388)
		sig_ram_VERS(4)
		sig_fnc_OWN(474)
		sig_ram_APP(5)
		sig_fnc_DATE(99)
		sig_ram_MKTA(4)
		sig_ram_MKTB(3)
		sig_ram_CABIN(7)
		sig_ram_BKG(6);
sig_rule(0000080) <= 
		sig_fnc_RTD(1029)
		sig_ram_VERS(0)
		sig_fnc_OWN(948)
		sig_ram_APP(4)
		sig_fnc_DATE(86)
		sig_ram_MKTA(30)
		sig_ram_MKTB(4)
		sig_ram_CABIN(6)
		sig_ram_BKG(16);
sig_rule(0000081) <= 
		sig_fnc_RTD(1814)
		sig_ram_VERS(1)
		sig_fnc_OWN(555)
		sig_ram_APP(43)
		sig_fnc_DATE(92)
		sig_ram_MKTA(25)
		sig_ram_MKTB(27)
		sig_ram_CABIN(4)
		sig_ram_BKG(7);
sig_rule(0000082) <= 
		sig_fnc_RTD(1786)
		sig_ram_VERS(3)
		sig_fnc_OWN(1029)
		sig_ram_APP(40)
		sig_fnc_DATE(76)
		sig_ram_MKTA(5)
		sig_ram_MKTB(6)
		sig_ram_CABIN(4)
		sig_ram_BKG(6);
sig_rule(0000083) <= 
		sig_fnc_RTD(35)
		sig_ram_VERS(2)
		sig_fnc_OWN(1003)
		sig_ram_APP(40)
		sig_fnc_DATE(11)
		sig_ram_MKTA(8)
		sig_ram_MKTB(2)
		sig_ram_CABIN(3)
		sig_ram_BKG(3);
sig_rule(0000084) <= 
		sig_fnc_RTD(2420)
		sig_ram_VERS(4)
		sig_fnc_OWN(1006)
		sig_ram_APP(33)
		sig_fnc_DATE(10)
		sig_ram_MKTA(21)
		sig_ram_MKTB(19)
		sig_ram_CABIN(1)
		sig_ram_BKG(9);
sig_rule(0000085) <= 
		sig_fnc_RTD(956)
		sig_ram_VERS(1)
		sig_fnc_OWN(544)
		sig_ram_APP(27)
		sig_fnc_DATE(70)
		sig_ram_MKTA(27)
		sig_ram_MKTB(16)
		sig_ram_CABIN(3)
		sig_ram_BKG(15);
sig_rule(0000086) <= 
		sig_fnc_RTD(147)
		sig_ram_VERS(0)
		sig_fnc_OWN(238)
		sig_ram_APP(8)
		sig_fnc_DATE(26)
		sig_ram_MKTA(20)
		sig_ram_MKTB(8)
		sig_ram_CABIN(7)
		sig_ram_BKG(18);
sig_rule(0000087) <= 
		sig_fnc_RTD(244)
		sig_ram_VERS(2)
		sig_fnc_OWN(567)
		sig_ram_APP(19)
		sig_fnc_DATE(50)
		sig_ram_MKTA(13)
		sig_ram_MKTB(21)
		sig_ram_CABIN(2)
		sig_ram_BKG(13);
sig_rule(0000088) <= 
		sig_fnc_RTD(527)
		sig_ram_VERS(3)
		sig_fnc_OWN(621)
		sig_ram_APP(8)
		sig_fnc_DATE(66)
		sig_ram_MKTA(6)
		sig_ram_MKTB(3)
		sig_ram_CABIN(5)
		sig_ram_BKG(18);
sig_rule(0000089) <= 
		sig_fnc_RTD(2115)
		sig_ram_VERS(1)
		sig_fnc_OWN(668)
		sig_ram_APP(24)
		sig_fnc_DATE(9)
		sig_ram_MKTA(8)
		sig_ram_MKTB(4)
		sig_ram_CABIN(1)
		sig_ram_BKG(14);
sig_rule(0000090) <= 
		sig_fnc_RTD(2765)
		sig_ram_VERS(2)
		sig_fnc_OWN(896)
		sig_ram_APP(20)
		sig_fnc_DATE(31)
		sig_ram_MKTA(5)
		sig_ram_MKTB(20)
		sig_ram_CABIN(1)
		sig_ram_BKG(9);
sig_rule(0000091) <= 
		sig_fnc_RTD(1013)
		sig_ram_VERS(1)
		sig_fnc_OWN(928)
		sig_ram_APP(19)
		sig_fnc_DATE(98)
		sig_ram_MKTA(19)
		sig_ram_MKTB(2)
		sig_ram_CABIN(7)
		sig_ram_BKG(24);
sig_rule(0000092) <= 
		sig_fnc_RTD(2148)
		sig_ram_VERS(1)
		sig_fnc_OWN(578)
		sig_ram_APP(34)
		sig_fnc_DATE(46)
		sig_ram_MKTA(23)
		sig_ram_MKTB(10)
		sig_ram_CABIN(4)
		sig_ram_BKG(7);
sig_rule(0000093) <= 
		sig_fnc_RTD(541)
		sig_ram_VERS(4)
		sig_fnc_OWN(887)
		sig_ram_APP(27)
		sig_fnc_DATE(92)
		sig_ram_MKTA(3)
		sig_ram_MKTB(28)
		sig_ram_CABIN(1)
		sig_ram_BKG(19);
sig_rule(0000094) <= 
		sig_fnc_RTD(1392)
		sig_ram_VERS(4)
		sig_fnc_OWN(989)
		sig_ram_APP(42)
		sig_fnc_DATE(81)
		sig_ram_MKTA(14)
		sig_ram_MKTB(12)
		sig_ram_CABIN(7)
		sig_ram_BKG(10);
sig_rule(0000095) <= 
		sig_fnc_RTD(2416)
		sig_ram_VERS(1)
		sig_fnc_OWN(180)
		sig_ram_APP(25)
		sig_fnc_DATE(43)
		sig_ram_MKTA(11)
		sig_ram_MKTB(22)
		sig_ram_CABIN(2)
		sig_ram_BKG(1);
sig_rule(0000096) <= 
		sig_fnc_RTD(2339)
		sig_ram_VERS(0)
		sig_fnc_OWN(593)
		sig_ram_APP(18)
		sig_fnc_DATE(46)
		sig_ram_MKTA(26)
		sig_ram_MKTB(23)
		sig_ram_CABIN(7)
		sig_ram_BKG(3);
sig_rule(0000097) <= 
		sig_fnc_RTD(786)
		sig_ram_VERS(4)
		sig_fnc_OWN(745)
		sig_ram_APP(43)
		sig_fnc_DATE(35)
		sig_ram_MKTA(21)
		sig_ram_MKTB(10)
		sig_ram_CABIN(1)
		sig_ram_BKG(13);
sig_rule(0000098) <= 
		sig_fnc_RTD(788)
		sig_ram_VERS(4)
		sig_fnc_OWN(899)
		sig_ram_APP(36)
		sig_fnc_DATE(50)
		sig_ram_MKTA(28)
		sig_ram_MKTB(29)
		sig_ram_CABIN(6)
		sig_ram_BKG(16);
sig_rule(0000099) <= 
		sig_fnc_RTD(2523)
		sig_ram_VERS(0)
		sig_fnc_OWN(340)
		sig_ram_APP(9)
		sig_fnc_DATE(94)
		sig_ram_MKTA(31)
		sig_ram_MKTB(28)
		sig_ram_CABIN(0);
