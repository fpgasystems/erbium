library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

package cfg_engines is

    constant THE_CFG_ENGINES_NUMBER       : integer :=  9; -- Number of engines per bitstream

end cfg_engines;

package body cfg_engines is

end cfg_engines;