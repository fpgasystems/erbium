
entity mct_wrapper 